module sid_mem16(
  input clk,
  input w_enable,
  input[12:0] address,
  input[15:0] data_in,
  output bit[15:0] data_out
);

(* no_rw_check *)
bit [15:0] m[8095:0];

always @(posedge clk) begin
  if (w_enable)
    m[address[12:0]] <= data_in;
  else
    data_out <= m[address[12:0]];
end

// cat Street_Fighter.cycles | nl -w1 -n ln -s " " -i2 -v1 | \
// nl -w1 -=16'h%04x;\nmn ln -s " " -i2 -v0 | \
// sed 's/\(.*\) \(.*\) \(.*\) \(.*\) \(.*\)/\1 \3 \2 \5 \4/g' | \
// tr '\n' ' ' | xargs -L1 printf "m[13'd%s]=16'h%04x;\nm[13'd%s]=16'h%02x%02x;\n" \
// > /tmp/mem.txt

initial begin
/*
    m[0] = 16'h0156;
    m[1] = 16'h0f18;
    m[2] = 16'h4d7e;
    m[3] = 16'h0018;
    m[7] = 3;
    m[15] = 4;
    m[31] = 5;
    m[63] = 6;
    m[127] = 7;
    m[255] = 8;
    m[511] = 9;
    m[1023] = 10;
    m[2047] = 11;
    m[4095] = 12;
    m[8191] = 13;
    m[16383] = 14;
    m[32767] = 15;
*/

m[13'd0]=16'h0156;
m[13'd1]=16'h0f18;
m[13'd2]=16'h4d7e;
m[13'd3]=16'h0018;
m[13'd4]=16'h000a;
m[13'd5]=16'h0017;
m[13'd6]=16'h000a;
m[13'd7]=16'h0016;
m[13'd8]=16'h000a;
m[13'd9]=16'h0015;
m[13'd10]=16'h000a;
m[13'd11]=16'h0014;
m[13'd12]=16'h000a;
m[13'd13]=16'h0013;
m[13'd14]=16'h000a;
m[13'd15]=16'h0012;
m[13'd16]=16'h000a;
m[13'd17]=16'h0011;
m[13'd18]=16'h000a;
m[13'd19]=16'h0010;
m[13'd20]=16'h000a;
m[13'd21]=16'h000f;
m[13'd22]=16'h000a;
m[13'd23]=16'h000e;
m[13'd24]=16'h000a;
m[13'd25]=16'h000d;
m[13'd26]=16'h000a;
m[13'd27]=16'h000c;
m[13'd28]=16'h000a;
m[13'd29]=16'h000b;
m[13'd30]=16'h000a;
m[13'd31]=16'h000a;
m[13'd32]=16'h000a;
m[13'd33]=16'h0009;
m[13'd34]=16'h000a;
m[13'd35]=16'h0008;
m[13'd36]=16'h000a;
m[13'd37]=16'h0007;
m[13'd38]=16'h000a;
m[13'd39]=16'h0006;
m[13'd40]=16'h000a;
m[13'd41]=16'h0005;
m[13'd42]=16'h000a;
m[13'd43]=16'h0004;
m[13'd44]=16'h000a;
m[13'd45]=16'h0003;
m[13'd46]=16'h000a;
m[13'd47]=16'h0002;
m[13'd48]=16'h000a;
m[13'd49]=16'h0001;
m[13'd50]=16'h000a;
m[13'd51]=16'h0000;
m[13'd52]=16'h0010;
m[13'd53]=16'h5f18;
m[13'd54]=16'h4af4;
m[13'd55]=16'h000f;
m[13'd56]=16'h0009;
m[13'd57]=16'h000e;
m[13'd58]=16'h001b;
m[13'd59]=16'h0010;
m[13'd60]=16'h0010;
m[13'd61]=16'h0011;
m[13'd62]=16'h0015;
m[13'd63]=16'h0013;
m[13'd64]=16'h0009;
m[13'd65]=16'h0014;
m[13'd66]=16'h0007;
m[13'd67]=16'h0012;
m[13'd68]=16'h0009;
m[13'd69]=16'h4012;
m[13'd70]=16'h016b;
m[13'd71]=16'h0008;
m[13'd72]=16'h0009;
m[13'd73]=16'h0007;
m[13'd74]=16'h001b;
m[13'd75]=16'h0009;
m[13'd76]=16'h0010;
m[13'd77]=16'h000a;
m[13'd78]=16'h0015;
m[13'd79]=16'h000c;
m[13'd80]=16'h0009;
m[13'd81]=16'h000d;
m[13'd82]=16'h0007;
m[13'd83]=16'h000b;
m[13'd84]=16'h0009;
m[13'd85]=16'h400b;
m[13'd86]=16'h020c;
m[13'd87]=16'h0301;
m[13'd88]=16'h0009;
m[13'd89]=16'h9b00;
m[13'd90]=16'h001b;
m[13'd91]=16'h4002;
m[13'd92]=16'h0010;
m[13'd93]=16'h0003;
m[13'd94]=16'h0016;
m[13'd95]=16'h0905;
m[13'd96]=16'h000a;
m[13'd97]=16'h0906;
m[13'd98]=16'h0007;
m[13'd99]=16'h0004;
m[13'd100]=16'h000a;
m[13'd101]=16'h4104;
m[13'd102]=16'h0095;
m[13'd103]=16'h0003;
m[13'd104]=16'h0009;
m[13'd105]=16'h5002;
m[13'd106]=16'h47db;
m[13'd107]=16'h0003;
m[13'd108]=16'h0009;
m[13'd109]=16'h6002;
m[13'd110]=16'h4cbd;
m[13'd111]=16'h0003;
m[13'd112]=16'h0009;
m[13'd113]=16'h7002;
m[13'd114]=16'h4cc0;
m[13'd115]=16'h0003;
m[13'd116]=16'h0009;
m[13'd117]=16'h8002;
m[13'd118]=16'h4cc0;
m[13'd119]=16'h0003;
m[13'd120]=16'h0009;
m[13'd121]=16'h9002;
m[13'd122]=16'h4cbd;
m[13'd123]=16'h0003;
m[13'd124]=16'h0009;
m[13'd125]=16'ha002;
m[13'd126]=16'h4c9d;
m[13'd127]=16'h4004;
m[13'd128]=16'h004e;
m[13'd129]=16'h0003;
m[13'd130]=16'h0009;
m[13'd131]=16'hb002;
m[13'd132]=16'h4c59;
m[13'd133]=16'h4004;
m[13'd134]=16'h004e;
m[13'd135]=16'h0003;
m[13'd136]=16'h0009;
m[13'd137]=16'hc002;
m[13'd138]=16'h4c70;
m[13'd139]=16'h4004;
m[13'd140]=16'h004e;
m[13'd141]=16'h0003;
m[13'd142]=16'h0009;
m[13'd143]=16'hd002;
m[13'd144]=16'h4c73;
m[13'd145]=16'h4004;
m[13'd146]=16'h004e;
m[13'd147]=16'h0003;
m[13'd148]=16'h0009;
m[13'd149]=16'he002;
m[13'd150]=16'h4c70;
m[13'd151]=16'h4004;
m[13'd152]=16'h004e;
m[13'd153]=16'h0003;
m[13'd154]=16'h0009;
m[13'd155]=16'hf002;
m[13'd156]=16'h4c70;
m[13'd157]=16'h4004;
m[13'd158]=16'h004e;
m[13'd159]=16'h0103;
m[13'd160]=16'h0009;
m[13'd161]=16'h0002;
m[13'd162]=16'h4cef;
m[13'd163]=16'h0301;
m[13'd164]=16'h0009;
m[13'd165]=16'h9b00;
m[13'd166]=16'h001b;
m[13'd167]=16'h4002;
m[13'd168]=16'h0010;
m[13'd169]=16'h0003;
m[13'd170]=16'h0016;
m[13'd171]=16'h0905;
m[13'd172]=16'h000a;
m[13'd173]=16'h0906;
m[13'd174]=16'h0007;
m[13'd175]=16'h0004;
m[13'd176]=16'h000a;
m[13'd177]=16'h4104;
m[13'd178]=16'h0095;
m[13'd179]=16'h0003;
m[13'd180]=16'h0009;
m[13'd181]=16'h5002;
m[13'd182]=16'h4b83;
m[13'd183]=16'h0003;
m[13'd184]=16'h0009;
m[13'd185]=16'h6002;
m[13'd186]=16'h4cc0;
m[13'd187]=16'h0003;
m[13'd188]=16'h0009;
m[13'd189]=16'h7002;
m[13'd190]=16'h4cbd;
m[13'd191]=16'h0003;
m[13'd192]=16'h0009;
m[13'd193]=16'h8002;
m[13'd194]=16'h4cc0;
m[13'd195]=16'h0003;
m[13'd196]=16'h0009;
m[13'd197]=16'h9002;
m[13'd198]=16'h4cc0;
m[13'd199]=16'h0003;
m[13'd200]=16'h0009;
m[13'd201]=16'ha002;
m[13'd202]=16'h4c9a;
m[13'd203]=16'h4004;
m[13'd204]=16'h004e;
m[13'd205]=16'h0003;
m[13'd206]=16'h0009;
m[13'd207]=16'hb002;
m[13'd208]=16'h4c59;
m[13'd209]=16'h4004;
m[13'd210]=16'h004e;
m[13'd211]=16'h0003;
m[13'd212]=16'h0009;
m[13'd213]=16'hc002;
m[13'd214]=16'h4c73;
m[13'd215]=16'h4004;
m[13'd216]=16'h004e;
m[13'd217]=16'h0003;
m[13'd218]=16'h0009;
m[13'd219]=16'hd002;
m[13'd220]=16'h4c70;
m[13'd221]=16'h4004;
m[13'd222]=16'h004e;
m[13'd223]=16'h0003;
m[13'd224]=16'h0009;
m[13'd225]=16'he002;
m[13'd226]=16'h4c70;
m[13'd227]=16'h4004;
m[13'd228]=16'h004e;
m[13'd229]=16'h0003;
m[13'd230]=16'h0009;
m[13'd231]=16'hf002;
m[13'd232]=16'h4c73;
m[13'd233]=16'h4004;
m[13'd234]=16'h004e;
m[13'd235]=16'h0103;
m[13'd236]=16'h0009;
m[13'd237]=16'h0002;
m[13'd238]=16'h4cf9;
m[13'd239]=16'h0301;
m[13'd240]=16'h0009;
m[13'd241]=16'h9b00;
m[13'd242]=16'h001b;
m[13'd243]=16'h4002;
m[13'd244]=16'h0010;
m[13'd245]=16'h0003;
m[13'd246]=16'h0016;
m[13'd247]=16'h0905;
m[13'd248]=16'h000a;
m[13'd249]=16'h0906;
m[13'd250]=16'h0007;
m[13'd251]=16'h0004;
m[13'd252]=16'h000a;
m[13'd253]=16'h4104;
m[13'd254]=16'h008d;
m[13'd255]=16'h0003;
m[13'd256]=16'h0009;
m[13'd257]=16'h5002;
m[13'd258]=16'h4b78;
m[13'd259]=16'h0003;
m[13'd260]=16'h0009;
m[13'd261]=16'h6002;
m[13'd262]=16'h4cbe;
m[13'd263]=16'h0003;
m[13'd264]=16'h0009;
m[13'd265]=16'h7002;
m[13'd266]=16'h4cbe;
m[13'd267]=16'h0003;
m[13'd268]=16'h0009;
m[13'd269]=16'h8002;
m[13'd270]=16'h4cc1;
m[13'd271]=16'h0003;
m[13'd272]=16'h0009;
m[13'd273]=16'h9002;
m[13'd274]=16'h4cbe;
m[13'd275]=16'h0003;
m[13'd276]=16'h0009;
m[13'd277]=16'ha002;
m[13'd278]=16'h4d07;
m[13'd279]=16'h0401;
m[13'd280]=16'h0009;
m[13'd281]=16'h4900;
m[13'd282]=16'h001b;
m[13'd283]=16'h4002;
m[13'd284]=16'h0010;
m[13'd285]=16'h0003;
m[13'd286]=16'h0016;
m[13'd287]=16'h0905;
m[13'd288]=16'h000a;
m[13'd289]=16'h0906;
m[13'd290]=16'h0007;
m[13'd291]=16'h0004;
m[13'd292]=16'h000a;
m[13'd293]=16'h4104;
m[13'd294]=16'h008d;
m[13'd295]=16'h0003;
m[13'd296]=16'h0009;
m[13'd297]=16'h5002;
m[13'd298]=16'h4b84;
m[13'd299]=16'h0003;
m[13'd300]=16'h0009;
m[13'd301]=16'h6002;
m[13'd302]=16'h4cc1;
m[13'd303]=16'h0003;
m[13'd304]=16'h0009;
m[13'd305]=16'h7002;
m[13'd306]=16'h4cbe;
m[13'd307]=16'h0003;
m[13'd308]=16'h0009;
m[13'd309]=16'h8002;
m[13'd310]=16'h4cbe;
m[13'd311]=16'h0003;
m[13'd312]=16'h0009;
m[13'd313]=16'h9002;
m[13'd314]=16'h4cc1;
m[13'd315]=16'h0003;
m[13'd316]=16'h0009;
m[13'd317]=16'ha002;
m[13'd318]=16'h4d14;
m[13'd319]=16'h0301;
m[13'd320]=16'h0009;
m[13'd321]=16'h9b00;
m[13'd322]=16'h001b;
m[13'd323]=16'h4002;
m[13'd324]=16'h0010;
m[13'd325]=16'h0003;
m[13'd326]=16'h0016;
m[13'd327]=16'h0905;
m[13'd328]=16'h000a;
m[13'd329]=16'h0906;
m[13'd330]=16'h0007;
m[13'd331]=16'h0004;
m[13'd332]=16'h000a;
m[13'd333]=16'h4104;
m[13'd334]=16'h0095;
m[13'd335]=16'h0003;
m[13'd336]=16'h0009;
m[13'd337]=16'h5002;
m[13'd338]=16'h4b77;
m[13'd339]=16'h0003;
m[13'd340]=16'h0009;
m[13'd341]=16'h6002;
m[13'd342]=16'h4cc0;
m[13'd343]=16'h0003;
m[13'd344]=16'h0009;
m[13'd345]=16'h7002;
m[13'd346]=16'h4cbd;
m[13'd347]=16'h0003;
m[13'd348]=16'h0009;
m[13'd349]=16'h8002;
m[13'd350]=16'h4cc0;
m[13'd351]=16'h0003;
m[13'd352]=16'h0009;
m[13'd353]=16'h9002;
m[13'd354]=16'h4cc0;
m[13'd355]=16'h0003;
m[13'd356]=16'h0009;
m[13'd357]=16'ha002;
m[13'd358]=16'h4c9a;
m[13'd359]=16'h4004;
m[13'd360]=16'h004e;
m[13'd361]=16'h0003;
m[13'd362]=16'h0009;
m[13'd363]=16'hb002;
m[13'd364]=16'h4c59;
m[13'd365]=16'h4004;
m[13'd366]=16'h004e;
m[13'd367]=16'h0003;
m[13'd368]=16'h0009;
m[13'd369]=16'hc002;
m[13'd370]=16'h4c73;
m[13'd371]=16'h4004;
m[13'd372]=16'h004e;
m[13'd373]=16'h0003;
m[13'd374]=16'h0009;
m[13'd375]=16'hd002;
m[13'd376]=16'h4c70;
m[13'd377]=16'h4004;
m[13'd378]=16'h004e;
m[13'd379]=16'h0003;
m[13'd380]=16'h0009;
m[13'd381]=16'he002;
m[13'd382]=16'h4c70;
m[13'd383]=16'h4004;
m[13'd384]=16'h004e;
m[13'd385]=16'h0003;
m[13'd386]=16'h0009;
m[13'd387]=16'hf002;
m[13'd388]=16'h4c73;
m[13'd389]=16'h4004;
m[13'd390]=16'h004e;
m[13'd391]=16'h0103;
m[13'd392]=16'h0009;
m[13'd393]=16'h0002;
m[13'd394]=16'h4cf9;
m[13'd395]=16'h0301;
m[13'd396]=16'h0009;
m[13'd397]=16'h9b00;
m[13'd398]=16'h001b;
m[13'd399]=16'h4002;
m[13'd400]=16'h0010;
m[13'd401]=16'h0003;
m[13'd402]=16'h0016;
m[13'd403]=16'h0905;
m[13'd404]=16'h000a;
m[13'd405]=16'h0906;
m[13'd406]=16'h0007;
m[13'd407]=16'h0004;
m[13'd408]=16'h000a;
m[13'd409]=16'h4104;
m[13'd410]=16'h008d;
m[13'd411]=16'h0003;
m[13'd412]=16'h0009;
m[13'd413]=16'h5002;
m[13'd414]=16'h4b78;
m[13'd415]=16'h0003;
m[13'd416]=16'h0009;
m[13'd417]=16'h6002;
m[13'd418]=16'h4cbe;
m[13'd419]=16'h0003;
m[13'd420]=16'h0009;
m[13'd421]=16'h7002;
m[13'd422]=16'h4cbe;
m[13'd423]=16'h0003;
m[13'd424]=16'h0009;
m[13'd425]=16'h8002;
m[13'd426]=16'h4cc1;
m[13'd427]=16'h0003;
m[13'd428]=16'h0009;
m[13'd429]=16'h9002;
m[13'd430]=16'h4cbe;
m[13'd431]=16'h0003;
m[13'd432]=16'h0009;
m[13'd433]=16'ha002;
m[13'd434]=16'h4d07;
m[13'd435]=16'h0401;
m[13'd436]=16'h0009;
m[13'd437]=16'hd000;
m[13'd438]=16'h001b;
m[13'd439]=16'h4002;
m[13'd440]=16'h0010;
m[13'd441]=16'h0003;
m[13'd442]=16'h0016;
m[13'd443]=16'h0905;
m[13'd444]=16'h000a;
m[13'd445]=16'h0906;
m[13'd446]=16'h0007;
m[13'd447]=16'h0004;
m[13'd448]=16'h000a;
m[13'd449]=16'h4104;
m[13'd450]=16'h008d;
m[13'd451]=16'h0003;
m[13'd452]=16'h0009;
m[13'd453]=16'h5002;
m[13'd454]=16'h4b84;
m[13'd455]=16'h0003;
m[13'd456]=16'h0009;
m[13'd457]=16'h6002;
m[13'd458]=16'h4cc1;
m[13'd459]=16'h0003;
m[13'd460]=16'h0009;
m[13'd461]=16'h7002;
m[13'd462]=16'h4cbe;
m[13'd463]=16'h0003;
m[13'd464]=16'h0009;
m[13'd465]=16'h8002;
m[13'd466]=16'h4cbe;
m[13'd467]=16'h0003;
m[13'd468]=16'h0009;
m[13'd469]=16'h9002;
m[13'd470]=16'h4cc1;
m[13'd471]=16'h0003;
m[13'd472]=16'h0009;
m[13'd473]=16'ha002;
m[13'd474]=16'h4d07;
m[13'd475]=16'h0301;
m[13'd476]=16'h0009;
m[13'd477]=16'h9b00;
m[13'd478]=16'h001b;
m[13'd479]=16'h4002;
m[13'd480]=16'h0010;
m[13'd481]=16'h0003;
m[13'd482]=16'h0016;
m[13'd483]=16'h0905;
m[13'd484]=16'h000a;
m[13'd485]=16'h0906;
m[13'd486]=16'h0007;
m[13'd487]=16'h0004;
m[13'd488]=16'h000a;
m[13'd489]=16'h4104;
m[13'd490]=16'h008d;
m[13'd491]=16'h0003;
m[13'd492]=16'h0009;
m[13'd493]=16'h5002;
m[13'd494]=16'h4b84;
m[13'd495]=16'h0003;
m[13'd496]=16'h0009;
m[13'd497]=16'h6002;
m[13'd498]=16'h4cbe;
m[13'd499]=16'h0003;
m[13'd500]=16'h0009;
m[13'd501]=16'h7002;
m[13'd502]=16'h4cc1;
m[13'd503]=16'h0003;
m[13'd504]=16'h0009;
m[13'd505]=16'h8002;
m[13'd506]=16'h4cbe;
m[13'd507]=16'h0003;
m[13'd508]=16'h0009;
m[13'd509]=16'h9002;
m[13'd510]=16'h4cbe;
m[13'd511]=16'h0003;
m[13'd512]=16'h0009;
m[13'd513]=16'ha002;
m[13'd514]=16'h4d0a;
m[13'd515]=16'h0301;
m[13'd516]=16'h0009;
m[13'd517]=16'h9b00;
m[13'd518]=16'h001b;
m[13'd519]=16'h4002;
m[13'd520]=16'h0010;
m[13'd521]=16'h0003;
m[13'd522]=16'h0016;
m[13'd523]=16'h0905;
m[13'd524]=16'h000a;
m[13'd525]=16'h0906;
m[13'd526]=16'h0007;
m[13'd527]=16'h0004;
m[13'd528]=16'h000a;
m[13'd529]=16'h4104;
m[13'd530]=16'h008d;
m[13'd531]=16'h0003;
m[13'd532]=16'h0009;
m[13'd533]=16'h5002;
m[13'd534]=16'h4b84;
m[13'd535]=16'h0003;
m[13'd536]=16'h0009;
m[13'd537]=16'h6002;
m[13'd538]=16'h4cbe;
m[13'd539]=16'h0003;
m[13'd540]=16'h0009;
m[13'd541]=16'h7002;
m[13'd542]=16'h4cbe;
m[13'd543]=16'h0003;
m[13'd544]=16'h0009;
m[13'd545]=16'h8002;
m[13'd546]=16'h4cc1;
m[13'd547]=16'h0003;
m[13'd548]=16'h0009;
m[13'd549]=16'h9002;
m[13'd550]=16'h4cbe;
m[13'd551]=16'h0003;
m[13'd552]=16'h0009;
m[13'd553]=16'ha002;
m[13'd554]=16'h4d07;
m[13'd555]=16'h0401;
m[13'd556]=16'h0009;
m[13'd557]=16'h4900;
m[13'd558]=16'h001b;
m[13'd559]=16'h4002;
m[13'd560]=16'h0010;
m[13'd561]=16'h0003;
m[13'd562]=16'h0016;
m[13'd563]=16'h0905;
m[13'd564]=16'h000a;
m[13'd565]=16'h0906;
m[13'd566]=16'h0007;
m[13'd567]=16'h0004;
m[13'd568]=16'h000a;
m[13'd569]=16'h4104;
m[13'd570]=16'h008d;
m[13'd571]=16'h0003;
m[13'd572]=16'h0009;
m[13'd573]=16'h5002;
m[13'd574]=16'h4b84;
m[13'd575]=16'h0003;
m[13'd576]=16'h0009;
m[13'd577]=16'h6002;
m[13'd578]=16'h4cc1;
m[13'd579]=16'h0003;
m[13'd580]=16'h0009;
m[13'd581]=16'h7002;
m[13'd582]=16'h4cbe;
m[13'd583]=16'h0003;
m[13'd584]=16'h0009;
m[13'd585]=16'h8002;
m[13'd586]=16'h4cbe;
m[13'd587]=16'h0003;
m[13'd588]=16'h0009;
m[13'd589]=16'h9002;
m[13'd590]=16'h4cc1;
m[13'd591]=16'h0003;
m[13'd592]=16'h0009;
m[13'd593]=16'ha002;
m[13'd594]=16'h4d14;
m[13'd595]=16'h0301;
m[13'd596]=16'h0009;
m[13'd597]=16'h9b00;
m[13'd598]=16'h001b;
m[13'd599]=16'h4002;
m[13'd600]=16'h0010;
m[13'd601]=16'h0003;
m[13'd602]=16'h0016;
m[13'd603]=16'h0905;
m[13'd604]=16'h000a;
m[13'd605]=16'h0906;
m[13'd606]=16'h0007;
m[13'd607]=16'h0004;
m[13'd608]=16'h000a;
m[13'd609]=16'h4104;
m[13'd610]=16'h0095;
m[13'd611]=16'h0003;
m[13'd612]=16'h0009;
m[13'd613]=16'h5002;
m[13'd614]=16'h4b77;
m[13'd615]=16'h0003;
m[13'd616]=16'h0009;
m[13'd617]=16'h6002;
m[13'd618]=16'h4cc0;
m[13'd619]=16'h0003;
m[13'd620]=16'h0009;
m[13'd621]=16'h7002;
m[13'd622]=16'h4cbd;
m[13'd623]=16'h0003;
m[13'd624]=16'h0009;
m[13'd625]=16'h8002;
m[13'd626]=16'h4cc0;
m[13'd627]=16'h0003;
m[13'd628]=16'h0009;
m[13'd629]=16'h9002;
m[13'd630]=16'h4cc0;
m[13'd631]=16'h0003;
m[13'd632]=16'h0009;
m[13'd633]=16'ha002;
m[13'd634]=16'h4c9a;
m[13'd635]=16'h4004;
m[13'd636]=16'h004e;
m[13'd637]=16'h0003;
m[13'd638]=16'h0009;
m[13'd639]=16'hb002;
m[13'd640]=16'h4c59;
m[13'd641]=16'h4004;
m[13'd642]=16'h004e;
m[13'd643]=16'h0003;
m[13'd644]=16'h0009;
m[13'd645]=16'hc002;
m[13'd646]=16'h4c73;
m[13'd647]=16'h4004;
m[13'd648]=16'h004e;
m[13'd649]=16'h0003;
m[13'd650]=16'h0009;
m[13'd651]=16'hd002;
m[13'd652]=16'h4c70;
m[13'd653]=16'h4004;
m[13'd654]=16'h004e;
m[13'd655]=16'h0003;
m[13'd656]=16'h0009;
m[13'd657]=16'he002;
m[13'd658]=16'h4c70;
m[13'd659]=16'h4004;
m[13'd660]=16'h004e;
m[13'd661]=16'h0003;
m[13'd662]=16'h0009;
m[13'd663]=16'hf002;
m[13'd664]=16'h4c73;
m[13'd665]=16'h4004;
m[13'd666]=16'h004e;
m[13'd667]=16'h0103;
m[13'd668]=16'h0009;
m[13'd669]=16'h0002;
m[13'd670]=16'h4cf9;
m[13'd671]=16'h0301;
m[13'd672]=16'h0009;
m[13'd673]=16'h3600;
m[13'd674]=16'h001b;
m[13'd675]=16'h4002;
m[13'd676]=16'h0010;
m[13'd677]=16'h0003;
m[13'd678]=16'h0016;
m[13'd679]=16'h0905;
m[13'd680]=16'h000a;
m[13'd681]=16'h0906;
m[13'd682]=16'h0007;
m[13'd683]=16'h0004;
m[13'd684]=16'h000a;
m[13'd685]=16'h4104;
m[13'd686]=16'h008d;
m[13'd687]=16'h0003;
m[13'd688]=16'h0009;
m[13'd689]=16'h5002;
m[13'd690]=16'h4b78;
m[13'd691]=16'h0003;
m[13'd692]=16'h0009;
m[13'd693]=16'h6002;
m[13'd694]=16'h4cbe;
m[13'd695]=16'h0003;
m[13'd696]=16'h0009;
m[13'd697]=16'h7002;
m[13'd698]=16'h4cbe;
m[13'd699]=16'h0003;
m[13'd700]=16'h0009;
m[13'd701]=16'h8002;
m[13'd702]=16'h4cc1;
m[13'd703]=16'h0003;
m[13'd704]=16'h0009;
m[13'd705]=16'h9002;
m[13'd706]=16'h4cbe;
m[13'd707]=16'h0003;
m[13'd708]=16'h0009;
m[13'd709]=16'ha002;
m[13'd710]=16'h4bb8;
m[13'd711]=16'h4012;
m[13'd712]=16'h0066;
m[13'd713]=16'h400b;
m[13'd714]=16'h011a;
m[13'd715]=16'h0301;
m[13'd716]=16'h0009;
m[13'd717]=16'h9b00;
m[13'd718]=16'h001b;
m[13'd719]=16'h4002;
m[13'd720]=16'h0010;
m[13'd721]=16'h0003;
m[13'd722]=16'h0016;
m[13'd723]=16'h0905;
m[13'd724]=16'h000a;
m[13'd725]=16'h0906;
m[13'd726]=16'h0007;
m[13'd727]=16'h0004;
m[13'd728]=16'h000a;
m[13'd729]=16'h4104;
m[13'd730]=16'h0095;
m[13'd731]=16'h0003;
m[13'd732]=16'h0009;
m[13'd733]=16'h5002;
m[13'd734]=16'h4a3d;
m[13'd735]=16'h4012;
m[13'd736]=16'h005e;
m[13'd737]=16'h400b;
m[13'd738]=16'h00dc;
m[13'd739]=16'h0003;
m[13'd740]=16'h0009;
m[13'd741]=16'h6002;
m[13'd742]=16'h4b86;
m[13'd743]=16'h4012;
m[13'd744]=16'h005e;
m[13'd745]=16'h400b;
m[13'd746]=16'h00dc;
m[13'd747]=16'h0003;
m[13'd748]=16'h0009;
m[13'd749]=16'h7002;
m[13'd750]=16'h4b86;
m[13'd751]=16'h4012;
m[13'd752]=16'h005e;
m[13'd753]=16'h400b;
m[13'd754]=16'h00dc;
m[13'd755]=16'h0003;
m[13'd756]=16'h0009;
m[13'd757]=16'h8002;
m[13'd758]=16'h4b83;
m[13'd759]=16'h4012;
m[13'd760]=16'h005e;
m[13'd761]=16'h400b;
m[13'd762]=16'h00dc;
m[13'd763]=16'h0003;
m[13'd764]=16'h0009;
m[13'd765]=16'h9002;
m[13'd766]=16'h4b86;
m[13'd767]=16'h4012;
m[13'd768]=16'h005e;
m[13'd769]=16'h400b;
m[13'd770]=16'h00dc;
m[13'd771]=16'h0003;
m[13'd772]=16'h0009;
m[13'd773]=16'ha002;
m[13'd774]=16'h4c79;
m[13'd775]=16'h4004;
m[13'd776]=16'h004e;
m[13'd777]=16'h0003;
m[13'd778]=16'h0009;
m[13'd779]=16'hb002;
m[13'd780]=16'h4c59;
m[13'd781]=16'h4004;
m[13'd782]=16'h004e;
m[13'd783]=16'h0003;
m[13'd784]=16'h0009;
m[13'd785]=16'hc002;
m[13'd786]=16'h4c70;
m[13'd787]=16'h4004;
m[13'd788]=16'h004e;
m[13'd789]=16'h0003;
m[13'd790]=16'h0009;
m[13'd791]=16'hd002;
m[13'd792]=16'h4c70;
m[13'd793]=16'h4004;
m[13'd794]=16'h004e;
m[13'd795]=16'h0003;
m[13'd796]=16'h0009;
m[13'd797]=16'he002;
m[13'd798]=16'h4c73;
m[13'd799]=16'h4004;
m[13'd800]=16'h004e;
m[13'd801]=16'h0003;
m[13'd802]=16'h0009;
m[13'd803]=16'hf002;
m[13'd804]=16'h4c70;
m[13'd805]=16'h4004;
m[13'd806]=16'h004e;
m[13'd807]=16'h0103;
m[13'd808]=16'h0009;
m[13'd809]=16'h0002;
m[13'd810]=16'h4cec;
m[13'd811]=16'h0301;
m[13'd812]=16'h0009;
m[13'd813]=16'h9b00;
m[13'd814]=16'h001b;
m[13'd815]=16'h4002;
m[13'd816]=16'h0010;
m[13'd817]=16'h0003;
m[13'd818]=16'h0016;
m[13'd819]=16'h0905;
m[13'd820]=16'h000a;
m[13'd821]=16'h0906;
m[13'd822]=16'h0007;
m[13'd823]=16'h0004;
m[13'd824]=16'h000a;
m[13'd825]=16'h4104;
m[13'd826]=16'h0095;
m[13'd827]=16'h0003;
m[13'd828]=16'h0009;
m[13'd829]=16'h5002;
m[13'd830]=16'h4b86;
m[13'd831]=16'h0003;
m[13'd832]=16'h0009;
m[13'd833]=16'h6002;
m[13'd834]=16'h4cbd;
m[13'd835]=16'h0003;
m[13'd836]=16'h0009;
m[13'd837]=16'h7002;
m[13'd838]=16'h4cc0;
m[13'd839]=16'h0003;
m[13'd840]=16'h0009;
m[13'd841]=16'h8002;
m[13'd842]=16'h4cc0;
m[13'd843]=16'h0003;
m[13'd844]=16'h0009;
m[13'd845]=16'h9002;
m[13'd846]=16'h4cbd;
m[13'd847]=16'h0003;
m[13'd848]=16'h0009;
m[13'd849]=16'ha002;
m[13'd850]=16'h4c9d;
m[13'd851]=16'h4004;
m[13'd852]=16'h004e;
m[13'd853]=16'h0003;
m[13'd854]=16'h0009;
m[13'd855]=16'hb002;
m[13'd856]=16'h4c59;
m[13'd857]=16'h4004;
m[13'd858]=16'h004e;
m[13'd859]=16'h0003;
m[13'd860]=16'h0009;
m[13'd861]=16'hc002;
m[13'd862]=16'h4c70;
m[13'd863]=16'h4004;
m[13'd864]=16'h004e;
m[13'd865]=16'h0003;
m[13'd866]=16'h0009;
m[13'd867]=16'hd002;
m[13'd868]=16'h4c73;
m[13'd869]=16'h4004;
m[13'd870]=16'h004e;
m[13'd871]=16'h0003;
m[13'd872]=16'h0009;
m[13'd873]=16'he002;
m[13'd874]=16'h4c70;
m[13'd875]=16'h4004;
m[13'd876]=16'h004e;
m[13'd877]=16'h0003;
m[13'd878]=16'h0009;
m[13'd879]=16'hf002;
m[13'd880]=16'h4c70;
m[13'd881]=16'h4004;
m[13'd882]=16'h004e;
m[13'd883]=16'h0103;
m[13'd884]=16'h0009;
m[13'd885]=16'h0002;
m[13'd886]=16'h4cfc;
m[13'd887]=16'h0301;
m[13'd888]=16'h0009;
m[13'd889]=16'h9b00;
m[13'd890]=16'h001b;
m[13'd891]=16'h4002;
m[13'd892]=16'h0010;
m[13'd893]=16'h0003;
m[13'd894]=16'h0016;
m[13'd895]=16'h0905;
m[13'd896]=16'h000a;
m[13'd897]=16'h0906;
m[13'd898]=16'h0007;
m[13'd899]=16'h0004;
m[13'd900]=16'h000a;
m[13'd901]=16'h4104;
m[13'd902]=16'h008d;
m[13'd903]=16'h0003;
m[13'd904]=16'h0009;
m[13'd905]=16'h5002;
m[13'd906]=16'h4b75;
m[13'd907]=16'h0003;
m[13'd908]=16'h0009;
m[13'd909]=16'h6002;
m[13'd910]=16'h4cc1;
m[13'd911]=16'h0003;
m[13'd912]=16'h0009;
m[13'd913]=16'h7002;
m[13'd914]=16'h4cbe;
m[13'd915]=16'h0003;
m[13'd916]=16'h0009;
m[13'd917]=16'h8002;
m[13'd918]=16'h4cbe;
m[13'd919]=16'h0003;
m[13'd920]=16'h0009;
m[13'd921]=16'h9002;
m[13'd922]=16'h4cc1;
m[13'd923]=16'h0003;
m[13'd924]=16'h0009;
m[13'd925]=16'ha002;
m[13'd926]=16'h4d07;
m[13'd927]=16'h0401;
m[13'd928]=16'h0009;
m[13'd929]=16'h4900;
m[13'd930]=16'h001b;
m[13'd931]=16'h4002;
m[13'd932]=16'h0010;
m[13'd933]=16'h0003;
m[13'd934]=16'h0016;
m[13'd935]=16'h0905;
m[13'd936]=16'h000a;
m[13'd937]=16'h0906;
m[13'd938]=16'h0007;
m[13'd939]=16'h0004;
m[13'd940]=16'h000a;
m[13'd941]=16'h4104;
m[13'd942]=16'h008d;
m[13'd943]=16'h0003;
m[13'd944]=16'h0009;
m[13'd945]=16'h5002;
m[13'd946]=16'h4b84;
m[13'd947]=16'h0003;
m[13'd948]=16'h0009;
m[13'd949]=16'h6002;
m[13'd950]=16'h4cbe;
m[13'd951]=16'h0003;
m[13'd952]=16'h0009;
m[13'd953]=16'h7002;
m[13'd954]=16'h4cc1;
m[13'd955]=16'h0003;
m[13'd956]=16'h0009;
m[13'd957]=16'h8002;
m[13'd958]=16'h4cbe;
m[13'd959]=16'h0003;
m[13'd960]=16'h0009;
m[13'd961]=16'h9002;
m[13'd962]=16'h4cbe;
m[13'd963]=16'h0003;
m[13'd964]=16'h0009;
m[13'd965]=16'ha002;
m[13'd966]=16'h4d17;
m[13'd967]=16'h0301;
m[13'd968]=16'h0009;
m[13'd969]=16'h9b00;
m[13'd970]=16'h001b;
m[13'd971]=16'h4002;
m[13'd972]=16'h0010;
m[13'd973]=16'h0003;
m[13'd974]=16'h0016;
m[13'd975]=16'h0905;
m[13'd976]=16'h000a;
m[13'd977]=16'h0906;
m[13'd978]=16'h0007;
m[13'd979]=16'h0004;
m[13'd980]=16'h000a;
m[13'd981]=16'h4104;
m[13'd982]=16'h0095;
m[13'd983]=16'h0003;
m[13'd984]=16'h0009;
m[13'd985]=16'h5002;
m[13'd986]=16'h4b77;
m[13'd987]=16'h0003;
m[13'd988]=16'h0009;
m[13'd989]=16'h6002;
m[13'd990]=16'h4cbd;
m[13'd991]=16'h0003;
m[13'd992]=16'h0009;
m[13'd993]=16'h7002;
m[13'd994]=16'h4cc0;
m[13'd995]=16'h0003;
m[13'd996]=16'h0009;
m[13'd997]=16'h8002;
m[13'd998]=16'h4cc0;
m[13'd999]=16'h0003;
m[13'd1000]=16'h0009;
m[13'd1001]=16'h9002;
m[13'd1002]=16'h4cbd;
m[13'd1003]=16'h0003;
m[13'd1004]=16'h0009;
m[13'd1005]=16'ha002;
m[13'd1006]=16'h4c9d;
m[13'd1007]=16'h4004;
m[13'd1008]=16'h004e;
m[13'd1009]=16'h0003;
m[13'd1010]=16'h0009;
m[13'd1011]=16'hb002;
m[13'd1012]=16'h4c59;
m[13'd1013]=16'h4004;
m[13'd1014]=16'h004e;
m[13'd1015]=16'h0003;
m[13'd1016]=16'h0009;
m[13'd1017]=16'hc002;
m[13'd1018]=16'h4c70;
m[13'd1019]=16'h4004;
m[13'd1020]=16'h004e;
m[13'd1021]=16'h0003;
m[13'd1022]=16'h0009;
m[13'd1023]=16'hd002;
m[13'd1024]=16'h4c73;
m[13'd1025]=16'h4004;
m[13'd1026]=16'h004e;
m[13'd1027]=16'h0003;
m[13'd1028]=16'h0009;
m[13'd1029]=16'he002;
m[13'd1030]=16'h4c70;
m[13'd1031]=16'h4004;
m[13'd1032]=16'h004e;
m[13'd1033]=16'h0003;
m[13'd1034]=16'h0009;
m[13'd1035]=16'hf002;
m[13'd1036]=16'h4c70;
m[13'd1037]=16'h4004;
m[13'd1038]=16'h004e;
m[13'd1039]=16'h0103;
m[13'd1040]=16'h0009;
m[13'd1041]=16'h0002;
m[13'd1042]=16'h4cfc;
m[13'd1043]=16'h0401;
m[13'd1044]=16'h0009;
m[13'd1045]=16'hd000;
m[13'd1046]=16'h001b;
m[13'd1047]=16'h4002;
m[13'd1048]=16'h0010;
m[13'd1049]=16'h0003;
m[13'd1050]=16'h0016;
m[13'd1051]=16'h0905;
m[13'd1052]=16'h000a;
m[13'd1053]=16'h0906;
m[13'd1054]=16'h0007;
m[13'd1055]=16'h0004;
m[13'd1056]=16'h000a;
m[13'd1057]=16'h4104;
m[13'd1058]=16'h008d;
m[13'd1059]=16'h0003;
m[13'd1060]=16'h0009;
m[13'd1061]=16'h5002;
m[13'd1062]=16'h4b75;
m[13'd1063]=16'h0003;
m[13'd1064]=16'h0009;
m[13'd1065]=16'h6002;
m[13'd1066]=16'h4cc1;
m[13'd1067]=16'h0003;
m[13'd1068]=16'h0009;
m[13'd1069]=16'h7002;
m[13'd1070]=16'h4cbe;
m[13'd1071]=16'h0003;
m[13'd1072]=16'h0009;
m[13'd1073]=16'h8002;
m[13'd1074]=16'h4cbe;
m[13'd1075]=16'h0003;
m[13'd1076]=16'h0009;
m[13'd1077]=16'h9002;
m[13'd1078]=16'h4cc1;
m[13'd1079]=16'h0003;
m[13'd1080]=16'h0009;
m[13'd1081]=16'ha002;
m[13'd1082]=16'h4d07;
m[13'd1083]=16'h0501;
m[13'd1084]=16'h0009;
m[13'd1085]=16'h1900;
m[13'd1086]=16'h001b;
m[13'd1087]=16'h4002;
m[13'd1088]=16'h0010;
m[13'd1089]=16'h0003;
m[13'd1090]=16'h0016;
m[13'd1091]=16'h0905;
m[13'd1092]=16'h000a;
m[13'd1093]=16'h0906;
m[13'd1094]=16'h0007;
m[13'd1095]=16'h0004;
m[13'd1096]=16'h000a;
m[13'd1097]=16'h4104;
m[13'd1098]=16'h008d;
m[13'd1099]=16'h0003;
m[13'd1100]=16'h0009;
m[13'd1101]=16'h5002;
m[13'd1102]=16'h4b84;
m[13'd1103]=16'h0003;
m[13'd1104]=16'h0009;
m[13'd1105]=16'h6002;
m[13'd1106]=16'h4cbe;
m[13'd1107]=16'h0003;
m[13'd1108]=16'h0009;
m[13'd1109]=16'h7002;
m[13'd1110]=16'h4cc1;
m[13'd1111]=16'h0003;
m[13'd1112]=16'h0009;
m[13'd1113]=16'h8002;
m[13'd1114]=16'h4cbe;
m[13'd1115]=16'h0003;
m[13'd1116]=16'h0009;
m[13'd1117]=16'h9002;
m[13'd1118]=16'h4cbe;
m[13'd1119]=16'h0003;
m[13'd1120]=16'h0009;
m[13'd1121]=16'ha002;
m[13'd1122]=16'h4d0a;
m[13'd1123]=16'h0501;
m[13'd1124]=16'h0009;
m[13'd1125]=16'h6700;
m[13'd1126]=16'h001b;
m[13'd1127]=16'h4002;
m[13'd1128]=16'h0010;
m[13'd1129]=16'h0003;
m[13'd1130]=16'h0016;
m[13'd1131]=16'h0905;
m[13'd1132]=16'h000a;
m[13'd1133]=16'h0906;
m[13'd1134]=16'h0007;
m[13'd1135]=16'h0004;
m[13'd1136]=16'h000a;
m[13'd1137]=16'h4104;
m[13'd1138]=16'h008d;
m[13'd1139]=16'h0003;
m[13'd1140]=16'h0009;
m[13'd1141]=16'h5002;
m[13'd1142]=16'h4b84;
m[13'd1143]=16'h0003;
m[13'd1144]=16'h0009;
m[13'd1145]=16'h6002;
m[13'd1146]=16'h4cbe;
m[13'd1147]=16'h0003;
m[13'd1148]=16'h0009;
m[13'd1149]=16'h7002;
m[13'd1150]=16'h4cbe;
m[13'd1151]=16'h0003;
m[13'd1152]=16'h0009;
m[13'd1153]=16'h8002;
m[13'd1154]=16'h4cc1;
m[13'd1155]=16'h0003;
m[13'd1156]=16'h0009;
m[13'd1157]=16'h9002;
m[13'd1158]=16'h4cbe;
m[13'd1159]=16'h0003;
m[13'd1160]=16'h0009;
m[13'd1161]=16'ha002;
m[13'd1162]=16'h4d15;
m[13'd1163]=16'h0601;
m[13'd1164]=16'h0009;
m[13'd1165]=16'h6c00;
m[13'd1166]=16'h001b;
m[13'd1167]=16'h4002;
m[13'd1168]=16'h0010;
m[13'd1169]=16'h0003;
m[13'd1170]=16'h0016;
m[13'd1171]=16'h0905;
m[13'd1172]=16'h000a;
m[13'd1173]=16'h0906;
m[13'd1174]=16'h0007;
m[13'd1175]=16'h0004;
m[13'd1176]=16'h000a;
m[13'd1177]=16'h4104;
m[13'd1178]=16'h0095;
m[13'd1179]=16'h0003;
m[13'd1180]=16'h0009;
m[13'd1181]=16'h5002;
m[13'd1182]=16'h4b77;
m[13'd1183]=16'h0003;
m[13'd1184]=16'h0009;
m[13'd1185]=16'h6002;
m[13'd1186]=16'h4cc0;
m[13'd1187]=16'h0003;
m[13'd1188]=16'h0009;
m[13'd1189]=16'h7002;
m[13'd1190]=16'h4cbd;
m[13'd1191]=16'h0003;
m[13'd1192]=16'h0009;
m[13'd1193]=16'h8002;
m[13'd1194]=16'h4cc0;
m[13'd1195]=16'h0003;
m[13'd1196]=16'h0009;
m[13'd1197]=16'h9002;
m[13'd1198]=16'h4cc0;
m[13'd1199]=16'h0003;
m[13'd1200]=16'h0009;
m[13'd1201]=16'ha002;
m[13'd1202]=16'h4c9a;
m[13'd1203]=16'h4004;
m[13'd1204]=16'h004e;
m[13'd1205]=16'h0003;
m[13'd1206]=16'h0009;
m[13'd1207]=16'hb002;
m[13'd1208]=16'h4c59;
m[13'd1209]=16'h4004;
m[13'd1210]=16'h004e;
m[13'd1211]=16'h0003;
m[13'd1212]=16'h0009;
m[13'd1213]=16'hc002;
m[13'd1214]=16'h4c73;
m[13'd1215]=16'h4004;
m[13'd1216]=16'h004e;
m[13'd1217]=16'h0003;
m[13'd1218]=16'h0009;
m[13'd1219]=16'hd002;
m[13'd1220]=16'h4c70;
m[13'd1221]=16'h4004;
m[13'd1222]=16'h004e;
m[13'd1223]=16'h0003;
m[13'd1224]=16'h0009;
m[13'd1225]=16'he002;
m[13'd1226]=16'h4c70;
m[13'd1227]=16'h4004;
m[13'd1228]=16'h004e;
m[13'd1229]=16'h0003;
m[13'd1230]=16'h0009;
m[13'd1231]=16'hf002;
m[13'd1232]=16'h4c73;
m[13'd1233]=16'h4004;
m[13'd1234]=16'h004e;
m[13'd1235]=16'h0103;
m[13'd1236]=16'h0009;
m[13'd1237]=16'h0002;
m[13'd1238]=16'h4cfa;
m[13'd1239]=16'h0501;
m[13'd1240]=16'h0009;
m[13'd1241]=16'hb900;
m[13'd1242]=16'h001b;
m[13'd1243]=16'h4002;
m[13'd1244]=16'h0010;
m[13'd1245]=16'h0003;
m[13'd1246]=16'h0016;
m[13'd1247]=16'h0905;
m[13'd1248]=16'h000a;
m[13'd1249]=16'h0906;
m[13'd1250]=16'h0007;
m[13'd1251]=16'h0004;
m[13'd1252]=16'h000a;
m[13'd1253]=16'h4104;
m[13'd1254]=16'h008d;
m[13'd1255]=16'h0003;
m[13'd1256]=16'h0009;
m[13'd1257]=16'h5002;
m[13'd1258]=16'h4b75;
m[13'd1259]=16'h0003;
m[13'd1260]=16'h0009;
m[13'd1261]=16'h6002;
m[13'd1262]=16'h4cc1;
m[13'd1263]=16'h0003;
m[13'd1264]=16'h0009;
m[13'd1265]=16'h7002;
m[13'd1266]=16'h4cbe;
m[13'd1267]=16'h0003;
m[13'd1268]=16'h0009;
m[13'd1269]=16'h8002;
m[13'd1270]=16'h4cbe;
m[13'd1271]=16'h0003;
m[13'd1272]=16'h0009;
m[13'd1273]=16'h9002;
m[13'd1274]=16'h4cc1;
m[13'd1275]=16'h0003;
m[13'd1276]=16'h0009;
m[13'd1277]=16'ha002;
m[13'd1278]=16'h4d08;
m[13'd1279]=16'h0601;
m[13'd1280]=16'h0009;
m[13'd1281]=16'h6c00;
m[13'd1282]=16'h001b;
m[13'd1283]=16'h4002;
m[13'd1284]=16'h0010;
m[13'd1285]=16'h0003;
m[13'd1286]=16'h0016;
m[13'd1287]=16'h0905;
m[13'd1288]=16'h000a;
m[13'd1289]=16'h0906;
m[13'd1290]=16'h0007;
m[13'd1291]=16'h0004;
m[13'd1292]=16'h000a;
m[13'd1293]=16'h4104;
m[13'd1294]=16'h008d;
m[13'd1295]=16'h0003;
m[13'd1296]=16'h0009;
m[13'd1297]=16'h5002;
m[13'd1298]=16'h4b84;
m[13'd1299]=16'h0003;
m[13'd1300]=16'h0009;
m[13'd1301]=16'h6002;
m[13'd1302]=16'h4cbe;
m[13'd1303]=16'h0003;
m[13'd1304]=16'h0009;
m[13'd1305]=16'h7002;
m[13'd1306]=16'h4cbe;
m[13'd1307]=16'h0003;
m[13'd1308]=16'h0009;
m[13'd1309]=16'h8002;
m[13'd1310]=16'h4cc1;
m[13'd1311]=16'h0003;
m[13'd1312]=16'h0009;
m[13'd1313]=16'h9002;
m[13'd1314]=16'h4cbe;
m[13'd1315]=16'h0003;
m[13'd1316]=16'h0009;
m[13'd1317]=16'ha002;
m[13'd1318]=16'h4d08;
m[13'd1319]=16'h0601;
m[13'd1320]=16'h0009;
m[13'd1321]=16'hce00;
m[13'd1322]=16'h001b;
m[13'd1323]=16'h4002;
m[13'd1324]=16'h0010;
m[13'd1325]=16'h0003;
m[13'd1326]=16'h0016;
m[13'd1327]=16'h0905;
m[13'd1328]=16'h000a;
m[13'd1329]=16'h0906;
m[13'd1330]=16'h0007;
m[13'd1331]=16'h0004;
m[13'd1332]=16'h000a;
m[13'd1333]=16'h4104;
m[13'd1334]=16'h008d;
m[13'd1335]=16'h0003;
m[13'd1336]=16'h0009;
m[13'd1337]=16'h5002;
m[13'd1338]=16'h4b84;
m[13'd1339]=16'h0003;
m[13'd1340]=16'h0009;
m[13'd1341]=16'h6002;
m[13'd1342]=16'h4cbe;
m[13'd1343]=16'h0003;
m[13'd1344]=16'h0009;
m[13'd1345]=16'h7002;
m[13'd1346]=16'h4cc1;
m[13'd1347]=16'h0003;
m[13'd1348]=16'h0009;
m[13'd1349]=16'h8002;
m[13'd1350]=16'h4cbe;
m[13'd1351]=16'h0003;
m[13'd1352]=16'h0009;
m[13'd1353]=16'h9002;
m[13'd1354]=16'h4cbe;
m[13'd1355]=16'h0003;
m[13'd1356]=16'h0009;
m[13'd1357]=16'ha002;
m[13'd1358]=16'h4ce0;
m[13'd1359]=16'h000f;
m[13'd1360]=16'h0009;
m[13'd1361]=16'h000e;
m[13'd1362]=16'h001b;
m[13'd1363]=16'h0010;
m[13'd1364]=16'h0010;
m[13'd1365]=16'h0011;
m[13'd1366]=16'h0015;
m[13'd1367]=16'h0013;
m[13'd1368]=16'h0009;
m[13'd1369]=16'h0014;
m[13'd1370]=16'h0007;
m[13'd1371]=16'h0012;
m[13'd1372]=16'h0009;
m[13'd1373]=16'h4012;
m[13'd1374]=16'h01c7;
m[13'd1375]=16'h0008;
m[13'd1376]=16'h0009;
m[13'd1377]=16'h0007;
m[13'd1378]=16'h001b;
m[13'd1379]=16'h0009;
m[13'd1380]=16'h0010;
m[13'd1381]=16'h000a;
m[13'd1382]=16'h0015;
m[13'd1383]=16'h000c;
m[13'd1384]=16'h0009;
m[13'd1385]=16'h000d;
m[13'd1386]=16'h0007;
m[13'd1387]=16'h000b;
m[13'd1388]=16'h0009;
m[13'd1389]=16'h400b;
m[13'd1390]=16'h0273;
m[13'd1391]=16'h0301;
m[13'd1392]=16'h0009;
m[13'd1393]=16'h9b00;
m[13'd1394]=16'h001b;
m[13'd1395]=16'h4002;
m[13'd1396]=16'h0010;
m[13'd1397]=16'h0003;
m[13'd1398]=16'h0016;
m[13'd1399]=16'h0905;
m[13'd1400]=16'h000a;
m[13'd1401]=16'h1906; // 0906
m[13'd1402]=16'h0007;
m[13'd1403]=16'h0004;
m[13'd1404]=16'h000a;
m[13'd1405]=16'h4104;
m[13'd1406]=16'h0095;
m[13'd1407]=16'h0003;
m[13'd1408]=16'h0009;
m[13'd1409]=16'h5002;
m[13'd1410]=16'h4633;
m[13'd1411]=16'h0000; // 4801
m[13'd1412]=16'h0007;
m[13'd1413]=16'h1801; // 0000
m[13'd1414]=16'h000e;
m[13'd1415]=16'h8104;
m[13'd1416]=16'h0060;
m[13'd1417]=16'h0003;
m[13'd1418]=16'h0009;
m[13'd1419]=16'h6002;
m[13'd1420]=16'h4c68;
m[13'd1421]=16'h0301;
m[13'd1422]=16'h0009;
m[13'd1423]=16'h9b00;
m[13'd1424]=16'h0018;
m[13'd1425]=16'h4104;
m[13'd1426]=16'h0060;
m[13'd1427]=16'h0003;
m[13'd1428]=16'h0009;
m[13'd1429]=16'h7002;
m[13'd1430]=16'h4c3e;
m[13'd1431]=16'h0301;
m[13'd1432]=16'h0009;
m[13'd1433]=16'h9b00;
m[13'd1434]=16'h0018;
m[13'd1435]=16'h4104;
m[13'd1436]=16'h0060;
m[13'd1437]=16'h0003;
m[13'd1438]=16'h0009;
m[13'd1439]=16'h8002;
m[13'd1440]=16'h4c3e;
m[13'd1441]=16'h0301;
m[13'd1442]=16'h0009;
m[13'd1443]=16'h9b00;
m[13'd1444]=16'h0018;
m[13'd1445]=16'h4104;
m[13'd1446]=16'h0060;
m[13'd1447]=16'h0003;
m[13'd1448]=16'h0009;
m[13'd1449]=16'h9002;
m[13'd1450]=16'h4c3e;
m[13'd1451]=16'h0301;
m[13'd1452]=16'h0009;
m[13'd1453]=16'h9b00;
m[13'd1454]=16'h0018;
m[13'd1455]=16'h4104;
m[13'd1456]=16'h0060;
m[13'd1457]=16'h0003;
m[13'd1458]=16'h0009;
m[13'd1459]=16'ha002;
m[13'd1460]=16'h4c56;
m[13'd1461]=16'h0301;
m[13'd1462]=16'h0009;
m[13'd1463]=16'h9b00;
m[13'd1464]=16'h0018;
m[13'd1465]=16'h4104;
m[13'd1466]=16'h0025;
m[13'd1467]=16'h4004;
m[13'd1468]=16'h004e;
m[13'd1469]=16'h0003;
m[13'd1470]=16'h0009;
m[13'd1471]=16'hb002;
m[13'd1472]=16'h4c12;
m[13'd1473]=16'h0301;
m[13'd1474]=16'h0009;
m[13'd1475]=16'h9b00;
m[13'd1476]=16'h0018;
m[13'd1477]=16'h4104;
m[13'd1478]=16'h0025;
m[13'd1479]=16'h4004;
m[13'd1480]=16'h004e;
m[13'd1481]=16'h0003;
m[13'd1482]=16'h0009;
m[13'd1483]=16'hc002;
m[13'd1484]=16'h4c2c;
m[13'd1485]=16'h0301;
m[13'd1486]=16'h0009;
m[13'd1487]=16'h9b00;
m[13'd1488]=16'h0018;
m[13'd1489]=16'h4104;
m[13'd1490]=16'h0025;
m[13'd1491]=16'h4004;
m[13'd1492]=16'h004e;
m[13'd1493]=16'h0003;
m[13'd1494]=16'h0009;
m[13'd1495]=16'hd002;
m[13'd1496]=16'h4c2c;
m[13'd1497]=16'h0301;
m[13'd1498]=16'h0009;
m[13'd1499]=16'h9b00;
m[13'd1500]=16'h0018;
m[13'd1501]=16'h4104;
m[13'd1502]=16'h0025;
m[13'd1503]=16'h4004;
m[13'd1504]=16'h004e;
m[13'd1505]=16'h0003;
m[13'd1506]=16'h0009;
m[13'd1507]=16'he002;
m[13'd1508]=16'h4c29;
m[13'd1509]=16'h0301;
m[13'd1510]=16'h0009;
m[13'd1511]=16'h9b00;
m[13'd1512]=16'h0018;
m[13'd1513]=16'h4104;
m[13'd1514]=16'h0025;
m[13'd1515]=16'h4004;
m[13'd1516]=16'h004e;
m[13'd1517]=16'h0003;
m[13'd1518]=16'h0009;
m[13'd1519]=16'hf002;
m[13'd1520]=16'h4c2c;
m[13'd1521]=16'h0301;
m[13'd1522]=16'h0009;
m[13'd1523]=16'h9b00;
m[13'd1524]=16'h0018;
m[13'd1525]=16'h4104;
m[13'd1526]=16'h0025;
m[13'd1527]=16'h4004;
m[13'd1528]=16'h004e;
m[13'd1529]=16'h0103;
m[13'd1530]=16'h0009;
m[13'd1531]=16'h0002;
m[13'd1532]=16'h4ccb;
m[13'd1533]=16'h0301;
m[13'd1534]=16'h0009;
m[13'd1535]=16'h9b00;
m[13'd1536]=16'h001b;
m[13'd1537]=16'h4002;
m[13'd1538]=16'h0010;
m[13'd1539]=16'h0003;
m[13'd1540]=16'h0016;
m[13'd1541]=16'h0905;
m[13'd1542]=16'h000a;
m[13'd1543]=16'h0906;
m[13'd1544]=16'h0007;
m[13'd1545]=16'h0004;
m[13'd1546]=16'h000a;
m[13'd1547]=16'h4104;
m[13'd1548]=16'h0095;
m[13'd1549]=16'h0003;
m[13'd1550]=16'h0009;
m[13'd1551]=16'h5002;
m[13'd1552]=16'h4b07;
m[13'd1553]=16'h4801;
m[13'd1554]=16'h0007;
m[13'd1555]=16'h0000;
m[13'd1556]=16'h000e;
m[13'd1557]=16'h8104;
m[13'd1558]=16'h0060;
m[13'd1559]=16'h0003;
m[13'd1560]=16'h0009;
m[13'd1561]=16'h6002;
m[13'd1562]=16'h4c68;
m[13'd1563]=16'h0301;
m[13'd1564]=16'h0009;
m[13'd1565]=16'h9b00;
m[13'd1566]=16'h0018;
m[13'd1567]=16'h4104;
m[13'd1568]=16'h0060;
m[13'd1569]=16'h0003;
m[13'd1570]=16'h0009;
m[13'd1571]=16'h7002;
m[13'd1572]=16'h4c3e;
m[13'd1573]=16'h0301;
m[13'd1574]=16'h0009;
m[13'd1575]=16'h9b00;
m[13'd1576]=16'h0018;
m[13'd1577]=16'h4104;
m[13'd1578]=16'h0060;
m[13'd1579]=16'h0003;
m[13'd1580]=16'h0009;
m[13'd1581]=16'h8002;
m[13'd1582]=16'h4c3e;
m[13'd1583]=16'h0301;
m[13'd1584]=16'h0009;
m[13'd1585]=16'h9b00;
m[13'd1586]=16'h0018;
m[13'd1587]=16'h4104;
m[13'd1588]=16'h0060;
m[13'd1589]=16'h0003;
m[13'd1590]=16'h0009;
m[13'd1591]=16'h9002;
m[13'd1592]=16'h4c3e;
m[13'd1593]=16'h0301;
m[13'd1594]=16'h0009;
m[13'd1595]=16'h9b00;
m[13'd1596]=16'h0018;
m[13'd1597]=16'h4104;
m[13'd1598]=16'h0060;
m[13'd1599]=16'h0003;
m[13'd1600]=16'h0009;
m[13'd1601]=16'ha002;
m[13'd1602]=16'h4c56;
m[13'd1603]=16'h0301;
m[13'd1604]=16'h0009;
m[13'd1605]=16'h9b00;
m[13'd1606]=16'h0018;
m[13'd1607]=16'h4104;
m[13'd1608]=16'h0025;
m[13'd1609]=16'h4004;
m[13'd1610]=16'h004e;
m[13'd1611]=16'h0003;
m[13'd1612]=16'h0009;
m[13'd1613]=16'hb002;
m[13'd1614]=16'h4c12;
m[13'd1615]=16'h0301;
m[13'd1616]=16'h0009;
m[13'd1617]=16'h9b00;
m[13'd1618]=16'h0018;
m[13'd1619]=16'h4104;
m[13'd1620]=16'h0025;
m[13'd1621]=16'h4004;
m[13'd1622]=16'h004e;
m[13'd1623]=16'h0003;
m[13'd1624]=16'h0009;
m[13'd1625]=16'hc002;
m[13'd1626]=16'h4c2c;
m[13'd1627]=16'h0301;
m[13'd1628]=16'h0009;
m[13'd1629]=16'h9b00;
m[13'd1630]=16'h0018;
m[13'd1631]=16'h4104;
m[13'd1632]=16'h0025;
m[13'd1633]=16'h4004;
m[13'd1634]=16'h004e;
m[13'd1635]=16'h0003;
m[13'd1636]=16'h0009;
m[13'd1637]=16'hd002;
m[13'd1638]=16'h4c2c;
m[13'd1639]=16'h0301;
m[13'd1640]=16'h0009;
m[13'd1641]=16'h9b00;
m[13'd1642]=16'h0018;
m[13'd1643]=16'h4104;
m[13'd1644]=16'h0025;
m[13'd1645]=16'h4004;
m[13'd1646]=16'h004e;
m[13'd1647]=16'h0003;
m[13'd1648]=16'h0009;
m[13'd1649]=16'he002;
m[13'd1650]=16'h4c29;
m[13'd1651]=16'h0301;
m[13'd1652]=16'h0009;
m[13'd1653]=16'h9b00;
m[13'd1654]=16'h0018;
m[13'd1655]=16'h4104;
m[13'd1656]=16'h0025;
m[13'd1657]=16'h4004;
m[13'd1658]=16'h004e;
m[13'd1659]=16'h0003;
m[13'd1660]=16'h0009;
m[13'd1661]=16'hf002;
m[13'd1662]=16'h4c2c;
m[13'd1663]=16'h0301;
m[13'd1664]=16'h0009;
m[13'd1665]=16'h9b00;
m[13'd1666]=16'h0018;
m[13'd1667]=16'h4104;
m[13'd1668]=16'h0025;
m[13'd1669]=16'h4004;
m[13'd1670]=16'h004e;
m[13'd1671]=16'h0103;
m[13'd1672]=16'h0009;
m[13'd1673]=16'h0002;
m[13'd1674]=16'h4cd8;
m[13'd1675]=16'h0301;
m[13'd1676]=16'h0009;
m[13'd1677]=16'h9b00;
m[13'd1678]=16'h001b;
m[13'd1679]=16'h4002;
m[13'd1680]=16'h0010;
m[13'd1681]=16'h0003;
m[13'd1682]=16'h0016;
m[13'd1683]=16'h0905;
m[13'd1684]=16'h000a;
m[13'd1685]=16'h0906;
m[13'd1686]=16'h0007;
m[13'd1687]=16'h0004;
m[13'd1688]=16'h000a;
m[13'd1689]=16'h4104;
m[13'd1690]=16'h008d;
m[13'd1691]=16'h0003;
m[13'd1692]=16'h0009;
m[13'd1693]=16'h5002;
m[13'd1694]=16'h4b01;
m[13'd1695]=16'h4801;
m[13'd1696]=16'h0007;
m[13'd1697]=16'h0000;
m[13'd1698]=16'h000e;
m[13'd1699]=16'h8104;
m[13'd1700]=16'h0058;
m[13'd1701]=16'h0003;
m[13'd1702]=16'h0009;
m[13'd1703]=16'h6002;
m[13'd1704]=16'h4c71;
m[13'd1705]=16'h0301;
m[13'd1706]=16'h0009;
m[13'd1707]=16'h9b00;
m[13'd1708]=16'h0018;
m[13'd1709]=16'h4104;
m[13'd1710]=16'h0058;
m[13'd1711]=16'h0003;
m[13'd1712]=16'h0009;
m[13'd1713]=16'h7002;
m[13'd1714]=16'h4c47;
m[13'd1715]=16'h0301;
m[13'd1716]=16'h0009;
m[13'd1717]=16'h9b00;
m[13'd1718]=16'h0018;
m[13'd1719]=16'h4104;
m[13'd1720]=16'h0058;
m[13'd1721]=16'h0003;
m[13'd1722]=16'h0009;
m[13'd1723]=16'h8002;
m[13'd1724]=16'h4c44;
m[13'd1725]=16'h0301;
m[13'd1726]=16'h0009;
m[13'd1727]=16'h9b00;
m[13'd1728]=16'h0018;
m[13'd1729]=16'h4104;
m[13'd1730]=16'h0058;
m[13'd1731]=16'h0003;
m[13'd1732]=16'h0009;
m[13'd1733]=16'h9002;
m[13'd1734]=16'h4c47;
m[13'd1735]=16'h0301;
m[13'd1736]=16'h0009;
m[13'd1737]=16'h9b00;
m[13'd1738]=16'h0018;
m[13'd1739]=16'h4104;
m[13'd1740]=16'h0058;
m[13'd1741]=16'h0003;
m[13'd1742]=16'h0009;
m[13'd1743]=16'ha002;
m[13'd1744]=16'h4ce6;
m[13'd1745]=16'h0401;
m[13'd1746]=16'h0009;
m[13'd1747]=16'h4900;
m[13'd1748]=16'h001b;
m[13'd1749]=16'h4002;
m[13'd1750]=16'h0010;
m[13'd1751]=16'h0003;
m[13'd1752]=16'h0016;
m[13'd1753]=16'h0905;
m[13'd1754]=16'h000a;
m[13'd1755]=16'h0906;
m[13'd1756]=16'h0007;
m[13'd1757]=16'h0004;
m[13'd1758]=16'h000a;
m[13'd1759]=16'h4104;
m[13'd1760]=16'h008d;
m[13'd1761]=16'h0003;
m[13'd1762]=16'h0009;
m[13'd1763]=16'h5002;
m[13'd1764]=16'h4b10;
m[13'd1765]=16'h4801;
m[13'd1766]=16'h0007;
m[13'd1767]=16'h0000;
m[13'd1768]=16'h000e;
m[13'd1769]=16'h8104;
m[13'd1770]=16'h0058;
m[13'd1771]=16'h0003;
m[13'd1772]=16'h0009;
m[13'd1773]=16'h6002;
m[13'd1774]=16'h4c6e;
m[13'd1775]=16'h0401;
m[13'd1776]=16'h0009;
m[13'd1777]=16'h4900;
m[13'd1778]=16'h0018;
m[13'd1779]=16'h4104;
m[13'd1780]=16'h0058;
m[13'd1781]=16'h0003;
m[13'd1782]=16'h0009;
m[13'd1783]=16'h7002;
m[13'd1784]=16'h4c47;
m[13'd1785]=16'h0401;
m[13'd1786]=16'h0009;
m[13'd1787]=16'h4900;
m[13'd1788]=16'h0018;
m[13'd1789]=16'h4104;
m[13'd1790]=16'h0058;
m[13'd1791]=16'h0003;
m[13'd1792]=16'h0009;
m[13'd1793]=16'h8002;
m[13'd1794]=16'h4c47;
m[13'd1795]=16'h0401;
m[13'd1796]=16'h0009;
m[13'd1797]=16'h4900;
m[13'd1798]=16'h0018;
m[13'd1799]=16'h4104;
m[13'd1800]=16'h0058;
m[13'd1801]=16'h0003;
m[13'd1802]=16'h0009;
m[13'd1803]=16'h9002;
m[13'd1804]=16'h4c44;
m[13'd1805]=16'h0401;
m[13'd1806]=16'h0009;
m[13'd1807]=16'h4900;
m[13'd1808]=16'h0018;
m[13'd1809]=16'h4104;
m[13'd1810]=16'h0058;
m[13'd1811]=16'h0003;
m[13'd1812]=16'h0009;
m[13'd1813]=16'ha002;
m[13'd1814]=16'h4cf3;
m[13'd1815]=16'h0301;
m[13'd1816]=16'h0009;
m[13'd1817]=16'h9b00;
m[13'd1818]=16'h001b;
m[13'd1819]=16'h4002;
m[13'd1820]=16'h0010;
m[13'd1821]=16'h0003;
m[13'd1822]=16'h0016;
m[13'd1823]=16'h0905;
m[13'd1824]=16'h000a;
m[13'd1825]=16'h0906;
m[13'd1826]=16'h0007;
m[13'd1827]=16'h0004;
m[13'd1828]=16'h000a;
m[13'd1829]=16'h4104;
m[13'd1830]=16'h0095;
m[13'd1831]=16'h0003;
m[13'd1832]=16'h0009;
m[13'd1833]=16'h5002;
m[13'd1834]=16'h4afb;
m[13'd1835]=16'h4801;
m[13'd1836]=16'h0007;
m[13'd1837]=16'h0000;
m[13'd1838]=16'h000e;
m[13'd1839]=16'h8104;
m[13'd1840]=16'h0060;
m[13'd1841]=16'h0003;
m[13'd1842]=16'h0009;
m[13'd1843]=16'h6002;
m[13'd1844]=16'h4c68;
m[13'd1845]=16'h0301;
m[13'd1846]=16'h0009;
m[13'd1847]=16'h9b00;
m[13'd1848]=16'h0018;
m[13'd1849]=16'h4104;
m[13'd1850]=16'h0060;
m[13'd1851]=16'h0003;
m[13'd1852]=16'h0009;
m[13'd1853]=16'h7002;
m[13'd1854]=16'h4c3e;
m[13'd1855]=16'h0301;
m[13'd1856]=16'h0009;
m[13'd1857]=16'h9b00;
m[13'd1858]=16'h0018;
m[13'd1859]=16'h4104;
m[13'd1860]=16'h0060;
m[13'd1861]=16'h0003;
m[13'd1862]=16'h0009;
m[13'd1863]=16'h8002;
m[13'd1864]=16'h4c3e;
m[13'd1865]=16'h0301;
m[13'd1866]=16'h0009;
m[13'd1867]=16'h9b00;
m[13'd1868]=16'h0018;
m[13'd1869]=16'h4104;
m[13'd1870]=16'h0060;
m[13'd1871]=16'h0003;
m[13'd1872]=16'h0009;
m[13'd1873]=16'h9002;
m[13'd1874]=16'h4c3e;
m[13'd1875]=16'h0301;
m[13'd1876]=16'h0009;
m[13'd1877]=16'h9b00;
m[13'd1878]=16'h0018;
m[13'd1879]=16'h4104;
m[13'd1880]=16'h0060;
m[13'd1881]=16'h0003;
m[13'd1882]=16'h0009;
m[13'd1883]=16'ha002;
m[13'd1884]=16'h4c56;
m[13'd1885]=16'h0301;
m[13'd1886]=16'h0009;
m[13'd1887]=16'h9b00;
m[13'd1888]=16'h0018;
m[13'd1889]=16'h4104;
m[13'd1890]=16'h0025;
m[13'd1891]=16'h4004;
m[13'd1892]=16'h004e;
m[13'd1893]=16'h0003;
m[13'd1894]=16'h0009;
m[13'd1895]=16'hb002;
m[13'd1896]=16'h4c12;
m[13'd1897]=16'h0301;
m[13'd1898]=16'h0009;
m[13'd1899]=16'h9b00;
m[13'd1900]=16'h0018;
m[13'd1901]=16'h4104;
m[13'd1902]=16'h0025;
m[13'd1903]=16'h4004;
m[13'd1904]=16'h004e;
m[13'd1905]=16'h0003;
m[13'd1906]=16'h0009;
m[13'd1907]=16'hc002;
m[13'd1908]=16'h4c2c;
m[13'd1909]=16'h0301;
m[13'd1910]=16'h0009;
m[13'd1911]=16'h9b00;
m[13'd1912]=16'h0018;
m[13'd1913]=16'h4104;
m[13'd1914]=16'h0025;
m[13'd1915]=16'h4004;
m[13'd1916]=16'h004e;
m[13'd1917]=16'h0003;
m[13'd1918]=16'h0009;
m[13'd1919]=16'hd002;
m[13'd1920]=16'h4c2c;
m[13'd1921]=16'h0301;
m[13'd1922]=16'h0009;
m[13'd1923]=16'h9b00;
m[13'd1924]=16'h0018;
m[13'd1925]=16'h4104;
m[13'd1926]=16'h0025;
m[13'd1927]=16'h4004;
m[13'd1928]=16'h004e;
m[13'd1929]=16'h0003;
m[13'd1930]=16'h0009;
m[13'd1931]=16'he002;
m[13'd1932]=16'h4c29;
m[13'd1933]=16'h0301;
m[13'd1934]=16'h0009;
m[13'd1935]=16'h9b00;
m[13'd1936]=16'h0018;
m[13'd1937]=16'h4104;
m[13'd1938]=16'h0025;
m[13'd1939]=16'h4004;
m[13'd1940]=16'h004e;
m[13'd1941]=16'h0003;
m[13'd1942]=16'h0009;
m[13'd1943]=16'hf002;
m[13'd1944]=16'h4c2c;
m[13'd1945]=16'h0301;
m[13'd1946]=16'h0009;
m[13'd1947]=16'h9b00;
m[13'd1948]=16'h0018;
m[13'd1949]=16'h4104;
m[13'd1950]=16'h0025;
m[13'd1951]=16'h4004;
m[13'd1952]=16'h004e;
m[13'd1953]=16'h0103;
m[13'd1954]=16'h0009;
m[13'd1955]=16'h0002;
m[13'd1956]=16'h4bd0;
m[13'd1957]=16'h400b;
m[13'd1958]=16'h011a;
m[13'd1959]=16'h0301;
m[13'd1960]=16'h0009;
m[13'd1961]=16'h9b00;
m[13'd1962]=16'h001b;
m[13'd1963]=16'h4002;
m[13'd1964]=16'h0010;
m[13'd1965]=16'h0003;
m[13'd1966]=16'h0016;
m[13'd1967]=16'h0905;
m[13'd1968]=16'h000a;
m[13'd1969]=16'h0906;
m[13'd1970]=16'h0007;
m[13'd1971]=16'h0004;
m[13'd1972]=16'h000a;
m[13'd1973]=16'h4104;
m[13'd1974]=16'h008d;
m[13'd1975]=16'h0003;
m[13'd1976]=16'h0009;
m[13'd1977]=16'h5002;
m[13'd1978]=16'h4aa1;
m[13'd1979]=16'h400b;
m[13'd1980]=16'h0060;
m[13'd1981]=16'h4801;
m[13'd1982]=16'h0007;
m[13'd1983]=16'h0000;
m[13'd1984]=16'h000e;
m[13'd1985]=16'h8104;
m[13'd1986]=16'h0058;
m[13'd1987]=16'h0003;
m[13'd1988]=16'h0009;
m[13'd1989]=16'h6002;
m[13'd1990]=16'h4bf3;
m[13'd1991]=16'h400b;
m[13'd1992]=16'h007e;
m[13'd1993]=16'h0301;
m[13'd1994]=16'h0009;
m[13'd1995]=16'h9b00;
m[13'd1996]=16'h0018;
m[13'd1997]=16'h4104;
m[13'd1998]=16'h0058;
m[13'd1999]=16'h0003;
m[13'd2000]=16'h0009;
m[13'd2001]=16'h7002;
m[13'd2002]=16'h4bc9;
m[13'd2003]=16'h400b;
m[13'd2004]=16'h007e;
m[13'd2005]=16'h0301;
m[13'd2006]=16'h0009;
m[13'd2007]=16'h9b00;
m[13'd2008]=16'h0018;
m[13'd2009]=16'h4104;
m[13'd2010]=16'h0058;
m[13'd2011]=16'h0003;
m[13'd2012]=16'h0009;
m[13'd2013]=16'h8002;
m[13'd2014]=16'h4bc6;
m[13'd2015]=16'h400b;
m[13'd2016]=16'h007e;
m[13'd2017]=16'h0301;
m[13'd2018]=16'h0009;
m[13'd2019]=16'h9b00;
m[13'd2020]=16'h0018;
m[13'd2021]=16'h4104;
m[13'd2022]=16'h0058;
m[13'd2023]=16'h0003;
m[13'd2024]=16'h0009;
m[13'd2025]=16'h9002;
m[13'd2026]=16'h4bc9;
m[13'd2027]=16'h400b;
m[13'd2028]=16'h007e;
m[13'd2029]=16'h0301;
m[13'd2030]=16'h0009;
m[13'd2031]=16'h9b00;
m[13'd2032]=16'h0018;
m[13'd2033]=16'h4104;
m[13'd2034]=16'h0058;
m[13'd2035]=16'h0003;
m[13'd2036]=16'h0009;
m[13'd2037]=16'ha002;
m[13'd2038]=16'h4cd4;
m[13'd2039]=16'h0401;
m[13'd2040]=16'h0009;
m[13'd2041]=16'hd000;
m[13'd2042]=16'h001b;
m[13'd2043]=16'h4002;
m[13'd2044]=16'h0010;
m[13'd2045]=16'h0003;
m[13'd2046]=16'h0016;
m[13'd2047]=16'h0905;
m[13'd2048]=16'h000a;
m[13'd2049]=16'h0906;
m[13'd2050]=16'h0007;
m[13'd2051]=16'h0004;
m[13'd2052]=16'h000a;
m[13'd2053]=16'h4104;
m[13'd2054]=16'h008d;
m[13'd2055]=16'h0003;
m[13'd2056]=16'h0009;
m[13'd2057]=16'h5002;
m[13'd2058]=16'h4b10;
m[13'd2059]=16'h4801;
m[13'd2060]=16'h0007;
m[13'd2061]=16'h0000;
m[13'd2062]=16'h000e;
m[13'd2063]=16'h8104;
m[13'd2064]=16'h0058;
m[13'd2065]=16'h0003;
m[13'd2066]=16'h0009;
m[13'd2067]=16'h6002;
m[13'd2068]=16'h4c6e;
m[13'd2069]=16'h0401;
m[13'd2070]=16'h0009;
m[13'd2071]=16'hd000;
m[13'd2072]=16'h0018;
m[13'd2073]=16'h4104;
m[13'd2074]=16'h0058;
m[13'd2075]=16'h0003;
m[13'd2076]=16'h0009;
m[13'd2077]=16'h7002;
m[13'd2078]=16'h4c47;
m[13'd2079]=16'h0401;
m[13'd2080]=16'h0009;
m[13'd2081]=16'hd000;
m[13'd2082]=16'h0018;
m[13'd2083]=16'h4104;
m[13'd2084]=16'h0058;
m[13'd2085]=16'h0003;
m[13'd2086]=16'h0009;
m[13'd2087]=16'h8002;
m[13'd2088]=16'h4c47;
m[13'd2089]=16'h0401;
m[13'd2090]=16'h0009;
m[13'd2091]=16'hd000;
m[13'd2092]=16'h0018;
m[13'd2093]=16'h4104;
m[13'd2094]=16'h0058;
m[13'd2095]=16'h0003;
m[13'd2096]=16'h0009;
m[13'd2097]=16'h9002;
m[13'd2098]=16'h4c44;
m[13'd2099]=16'h0401;
m[13'd2100]=16'h0009;
m[13'd2101]=16'hd000;
m[13'd2102]=16'h0018;
m[13'd2103]=16'h4104;
m[13'd2104]=16'h0058;
m[13'd2105]=16'h0003;
m[13'd2106]=16'h0009;
m[13'd2107]=16'ha002;
m[13'd2108]=16'h4ce6;
m[13'd2109]=16'h0301;
m[13'd2110]=16'h0009;
m[13'd2111]=16'h9b00;
m[13'd2112]=16'h001b;
m[13'd2113]=16'h4002;
m[13'd2114]=16'h0010;
m[13'd2115]=16'h0003;
m[13'd2116]=16'h0016;
m[13'd2117]=16'h0905;
m[13'd2118]=16'h000a;
m[13'd2119]=16'h0906;
m[13'd2120]=16'h0007;
m[13'd2121]=16'h0004;
m[13'd2122]=16'h000a;
m[13'd2123]=16'h4104;
m[13'd2124]=16'h008d;
m[13'd2125]=16'h0003;
m[13'd2126]=16'h0009;
m[13'd2127]=16'h5002;
m[13'd2128]=16'h4b10;
m[13'd2129]=16'h4801;
m[13'd2130]=16'h0007;
m[13'd2131]=16'h0000;
m[13'd2132]=16'h000e;
m[13'd2133]=16'h8104;
m[13'd2134]=16'h0058;
m[13'd2135]=16'h0003;
m[13'd2136]=16'h0009;
m[13'd2137]=16'h6002;
m[13'd2138]=16'h4c71;
m[13'd2139]=16'h0301;
m[13'd2140]=16'h0009;
m[13'd2141]=16'h9b00;
m[13'd2142]=16'h0018;
m[13'd2143]=16'h4104;
m[13'd2144]=16'h0058;
m[13'd2145]=16'h0003;
m[13'd2146]=16'h0009;
m[13'd2147]=16'h7002;
m[13'd2148]=16'h4c44;
m[13'd2149]=16'h0301;
m[13'd2150]=16'h0009;
m[13'd2151]=16'h9b00;
m[13'd2152]=16'h0018;
m[13'd2153]=16'h4104;
m[13'd2154]=16'h0058;
m[13'd2155]=16'h0003;
m[13'd2156]=16'h0009;
m[13'd2157]=16'h8002;
m[13'd2158]=16'h4c47;
m[13'd2159]=16'h0301;
m[13'd2160]=16'h0009;
m[13'd2161]=16'h9b00;
m[13'd2162]=16'h0018;
m[13'd2163]=16'h4104;
m[13'd2164]=16'h0058;
m[13'd2165]=16'h0003;
m[13'd2166]=16'h0009;
m[13'd2167]=16'h9002;
m[13'd2168]=16'h4c47;
m[13'd2169]=16'h0301;
m[13'd2170]=16'h0009;
m[13'd2171]=16'h9b00;
m[13'd2172]=16'h0018;
m[13'd2173]=16'h4104;
m[13'd2174]=16'h0058;
m[13'd2175]=16'h0003;
m[13'd2176]=16'h0009;
m[13'd2177]=16'ha002;
m[13'd2178]=16'h4ce3;
m[13'd2179]=16'h0301;
m[13'd2180]=16'h0009;
m[13'd2181]=16'h9b00;
m[13'd2182]=16'h001b;
m[13'd2183]=16'h4002;
m[13'd2184]=16'h0010;
m[13'd2185]=16'h0003;
m[13'd2186]=16'h0016;
m[13'd2187]=16'h0905;
m[13'd2188]=16'h000a;
m[13'd2189]=16'h0906;
m[13'd2190]=16'h0007;
m[13'd2191]=16'h0004;
m[13'd2192]=16'h000a;
m[13'd2193]=16'h4104;
m[13'd2194]=16'h008d;
m[13'd2195]=16'h0003;
m[13'd2196]=16'h0009;
m[13'd2197]=16'h5002;
m[13'd2198]=16'h4b10;
m[13'd2199]=16'h4801;
m[13'd2200]=16'h0007;
m[13'd2201]=16'h0000;
m[13'd2202]=16'h000e;
m[13'd2203]=16'h8104;
m[13'd2204]=16'h0058;
m[13'd2205]=16'h0003;
m[13'd2206]=16'h0009;
m[13'd2207]=16'h6002;
m[13'd2208]=16'h4c71;
m[13'd2209]=16'h0301;
m[13'd2210]=16'h0009;
m[13'd2211]=16'h9b00;
m[13'd2212]=16'h0018;
m[13'd2213]=16'h4104;
m[13'd2214]=16'h0058;
m[13'd2215]=16'h0003;
m[13'd2216]=16'h0009;
m[13'd2217]=16'h7002;
m[13'd2218]=16'h4c47;
m[13'd2219]=16'h0301;
m[13'd2220]=16'h0009;
m[13'd2221]=16'h9b00;
m[13'd2222]=16'h0018;
m[13'd2223]=16'h4104;
m[13'd2224]=16'h0058;
m[13'd2225]=16'h0003;
m[13'd2226]=16'h0009;
m[13'd2227]=16'h8002;
m[13'd2228]=16'h4c44;
m[13'd2229]=16'h0301;
m[13'd2230]=16'h0009;
m[13'd2231]=16'h9b00;
m[13'd2232]=16'h0018;
m[13'd2233]=16'h4104;
m[13'd2234]=16'h0058;
m[13'd2235]=16'h0003;
m[13'd2236]=16'h0009;
m[13'd2237]=16'h9002;
m[13'd2238]=16'h4c47;
m[13'd2239]=16'h0301;
m[13'd2240]=16'h0009;
m[13'd2241]=16'h9b00;
m[13'd2242]=16'h0018;
m[13'd2243]=16'h4104;
m[13'd2244]=16'h0058;
m[13'd2245]=16'h0003;
m[13'd2246]=16'h0009;
m[13'd2247]=16'ha002;
m[13'd2248]=16'h4ce6;
m[13'd2249]=16'h0401;
m[13'd2250]=16'h0009;
m[13'd2251]=16'h4900;
m[13'd2252]=16'h001b;
m[13'd2253]=16'h4002;
m[13'd2254]=16'h0010;
m[13'd2255]=16'h0003;
m[13'd2256]=16'h0016;
m[13'd2257]=16'h0905;
m[13'd2258]=16'h000a;
m[13'd2259]=16'h0906;
m[13'd2260]=16'h0007;
m[13'd2261]=16'h0004;
m[13'd2262]=16'h000a;
m[13'd2263]=16'h4104;
m[13'd2264]=16'h008d;
m[13'd2265]=16'h0003;
m[13'd2266]=16'h0009;
m[13'd2267]=16'h5002;
m[13'd2268]=16'h4b10;
m[13'd2269]=16'h4801;
m[13'd2270]=16'h0007;
m[13'd2271]=16'h0000;
m[13'd2272]=16'h000e;
m[13'd2273]=16'h8104;
m[13'd2274]=16'h0058;
m[13'd2275]=16'h0003;
m[13'd2276]=16'h0009;
m[13'd2277]=16'h6002;
m[13'd2278]=16'h4c6e;
m[13'd2279]=16'h0401;
m[13'd2280]=16'h0009;
m[13'd2281]=16'h4900;
m[13'd2282]=16'h0018;
m[13'd2283]=16'h4104;
m[13'd2284]=16'h0058;
m[13'd2285]=16'h0003;
m[13'd2286]=16'h0009;
m[13'd2287]=16'h7002;
m[13'd2288]=16'h4c47;
m[13'd2289]=16'h0401;
m[13'd2290]=16'h0009;
m[13'd2291]=16'h4900;
m[13'd2292]=16'h0018;
m[13'd2293]=16'h4104;
m[13'd2294]=16'h0058;
m[13'd2295]=16'h0003;
m[13'd2296]=16'h0009;
m[13'd2297]=16'h8002;
m[13'd2298]=16'h4c47;
m[13'd2299]=16'h0401;
m[13'd2300]=16'h0009;
m[13'd2301]=16'h4900;
m[13'd2302]=16'h0018;
m[13'd2303]=16'h4104;
m[13'd2304]=16'h0058;
m[13'd2305]=16'h0003;
m[13'd2306]=16'h0009;
m[13'd2307]=16'h9002;
m[13'd2308]=16'h4c44;
m[13'd2309]=16'h0401;
m[13'd2310]=16'h0009;
m[13'd2311]=16'h4900;
m[13'd2312]=16'h0018;
m[13'd2313]=16'h4104;
m[13'd2314]=16'h0058;
m[13'd2315]=16'h0003;
m[13'd2316]=16'h0009;
m[13'd2317]=16'ha002;
m[13'd2318]=16'h4cf3;
m[13'd2319]=16'h0301;
m[13'd2320]=16'h0009;
m[13'd2321]=16'h9b00;
m[13'd2322]=16'h001b;
m[13'd2323]=16'h4002;
m[13'd2324]=16'h0010;
m[13'd2325]=16'h0003;
m[13'd2326]=16'h0016;
m[13'd2327]=16'h0905;
m[13'd2328]=16'h000a;
m[13'd2329]=16'h0906;
m[13'd2330]=16'h0007;
m[13'd2331]=16'h0004;
m[13'd2332]=16'h000a;
m[13'd2333]=16'h4104;
m[13'd2334]=16'h0095;
m[13'd2335]=16'h0003;
m[13'd2336]=16'h0009;
m[13'd2337]=16'h5002;
m[13'd2338]=16'h4afb;
m[13'd2339]=16'h4801;
m[13'd2340]=16'h0007;
m[13'd2341]=16'h0000;
m[13'd2342]=16'h000e;
m[13'd2343]=16'h8104;
m[13'd2344]=16'h0060;
m[13'd2345]=16'h0003;
m[13'd2346]=16'h0009;
m[13'd2347]=16'h6002;
m[13'd2348]=16'h4c68;
m[13'd2349]=16'h0301;
m[13'd2350]=16'h0009;
m[13'd2351]=16'h9b00;
m[13'd2352]=16'h0018;
m[13'd2353]=16'h4104;
m[13'd2354]=16'h0060;
m[13'd2355]=16'h0003;
m[13'd2356]=16'h0009;
m[13'd2357]=16'h7002;
m[13'd2358]=16'h4c3e;
m[13'd2359]=16'h0301;
m[13'd2360]=16'h0009;
m[13'd2361]=16'h9b00;
m[13'd2362]=16'h0018;
m[13'd2363]=16'h4104;
m[13'd2364]=16'h0060;
m[13'd2365]=16'h0003;
m[13'd2366]=16'h0009;
m[13'd2367]=16'h8002;
m[13'd2368]=16'h4c3e;
m[13'd2369]=16'h0301;
m[13'd2370]=16'h0009;
m[13'd2371]=16'h9b00;
m[13'd2372]=16'h0018;
m[13'd2373]=16'h4104;
m[13'd2374]=16'h0060;
m[13'd2375]=16'h0003;
m[13'd2376]=16'h0009;
m[13'd2377]=16'h9002;
m[13'd2378]=16'h4c3e;
m[13'd2379]=16'h0301;
m[13'd2380]=16'h0009;
m[13'd2381]=16'h9b00;
m[13'd2382]=16'h0018;
m[13'd2383]=16'h4104;
m[13'd2384]=16'h0060;
m[13'd2385]=16'h0003;
m[13'd2386]=16'h0009;
m[13'd2387]=16'ha002;
m[13'd2388]=16'h4c56;
m[13'd2389]=16'h0301;
m[13'd2390]=16'h0009;
m[13'd2391]=16'h9b00;
m[13'd2392]=16'h0018;
m[13'd2393]=16'h4104;
m[13'd2394]=16'h0025;
m[13'd2395]=16'h4004;
m[13'd2396]=16'h004e;
m[13'd2397]=16'h0003;
m[13'd2398]=16'h0009;
m[13'd2399]=16'hb002;
m[13'd2400]=16'h4c12;
m[13'd2401]=16'h0301;
m[13'd2402]=16'h0009;
m[13'd2403]=16'h9b00;
m[13'd2404]=16'h0018;
m[13'd2405]=16'h4104;
m[13'd2406]=16'h0025;
m[13'd2407]=16'h4004;
m[13'd2408]=16'h004e;
m[13'd2409]=16'h0003;
m[13'd2410]=16'h0009;
m[13'd2411]=16'hc002;
m[13'd2412]=16'h4c2c;
m[13'd2413]=16'h0301;
m[13'd2414]=16'h0009;
m[13'd2415]=16'h9b00;
m[13'd2416]=16'h0018;
m[13'd2417]=16'h4104;
m[13'd2418]=16'h0025;
m[13'd2419]=16'h4004;
m[13'd2420]=16'h004e;
m[13'd2421]=16'h0003;
m[13'd2422]=16'h0009;
m[13'd2423]=16'hd002;
m[13'd2424]=16'h4c2c;
m[13'd2425]=16'h0301;
m[13'd2426]=16'h0009;
m[13'd2427]=16'h9b00;
m[13'd2428]=16'h0018;
m[13'd2429]=16'h4104;
m[13'd2430]=16'h0025;
m[13'd2431]=16'h4004;
m[13'd2432]=16'h004e;
m[13'd2433]=16'h0003;
m[13'd2434]=16'h0009;
m[13'd2435]=16'he002;
m[13'd2436]=16'h4c29;
m[13'd2437]=16'h0301;
m[13'd2438]=16'h0009;
m[13'd2439]=16'h9b00;
m[13'd2440]=16'h0018;
m[13'd2441]=16'h4104;
m[13'd2442]=16'h0025;
m[13'd2443]=16'h4004;
m[13'd2444]=16'h004e;
m[13'd2445]=16'h0003;
m[13'd2446]=16'h0009;
m[13'd2447]=16'hf002;
m[13'd2448]=16'h4c2c;
m[13'd2449]=16'h0301;
m[13'd2450]=16'h0009;
m[13'd2451]=16'h9b00;
m[13'd2452]=16'h0018;
m[13'd2453]=16'h4104;
m[13'd2454]=16'h0025;
m[13'd2455]=16'h4004;
m[13'd2456]=16'h004e;
m[13'd2457]=16'h0103;
m[13'd2458]=16'h0009;
m[13'd2459]=16'h0002;
m[13'd2460]=16'h4cd8;
m[13'd2461]=16'h0301;
m[13'd2462]=16'h0009;
m[13'd2463]=16'h3600;
m[13'd2464]=16'h001b;
m[13'd2465]=16'h4002;
m[13'd2466]=16'h0010;
m[13'd2467]=16'h0003;
m[13'd2468]=16'h0016;
m[13'd2469]=16'h0905;
m[13'd2470]=16'h000a;
m[13'd2471]=16'h0906;
m[13'd2472]=16'h0007;
m[13'd2473]=16'h0004;
m[13'd2474]=16'h000a;
m[13'd2475]=16'h4104;
m[13'd2476]=16'h008d;
m[13'd2477]=16'h0003;
m[13'd2478]=16'h0009;
m[13'd2479]=16'h5002;
m[13'd2480]=16'h4b01;
m[13'd2481]=16'h4801;
m[13'd2482]=16'h0007;
m[13'd2483]=16'h0000;
m[13'd2484]=16'h000e;
m[13'd2485]=16'h8104;
m[13'd2486]=16'h0058;
m[13'd2487]=16'h0003;
m[13'd2488]=16'h0009;
m[13'd2489]=16'h6002;
m[13'd2490]=16'h4c71;
m[13'd2491]=16'h0301;
m[13'd2492]=16'h0009;
m[13'd2493]=16'h3600;
m[13'd2494]=16'h0018;
m[13'd2495]=16'h4104;
m[13'd2496]=16'h0058;
m[13'd2497]=16'h0003;
m[13'd2498]=16'h0009;
m[13'd2499]=16'h7002;
m[13'd2500]=16'h4c47;
m[13'd2501]=16'h0301;
m[13'd2502]=16'h0009;
m[13'd2503]=16'h3600;
m[13'd2504]=16'h0018;
m[13'd2505]=16'h4104;
m[13'd2506]=16'h0058;
m[13'd2507]=16'h0003;
m[13'd2508]=16'h0009;
m[13'd2509]=16'h8002;
m[13'd2510]=16'h4c44;
m[13'd2511]=16'h0301;
m[13'd2512]=16'h0009;
m[13'd2513]=16'h3600;
m[13'd2514]=16'h0018;
m[13'd2515]=16'h4104;
m[13'd2516]=16'h0058;
m[13'd2517]=16'h0003;
m[13'd2518]=16'h0009;
m[13'd2519]=16'h9002;
m[13'd2520]=16'h4c47;
m[13'd2521]=16'h0301;
m[13'd2522]=16'h0009;
m[13'd2523]=16'h3600;
m[13'd2524]=16'h0018;
m[13'd2525]=16'h4104;
m[13'd2526]=16'h0058;
m[13'd2527]=16'h0003;
m[13'd2528]=16'h0009;
m[13'd2529]=16'ha002;
m[13'd2530]=16'h4b97;
m[13'd2531]=16'h4012;
m[13'd2532]=16'h012e;
m[13'd2533]=16'h0308;
m[13'd2534]=16'h0009;
m[13'd2535]=16'h6707;
m[13'd2536]=16'h001b;
m[13'd2537]=16'h8009;
m[13'd2538]=16'h0010;
m[13'd2539]=16'h000a;
m[13'd2540]=16'h0015;
m[13'd2541]=16'h090c;
m[13'd2542]=16'h0009;
m[13'd2543]=16'h080d;
m[13'd2544]=16'h0007;
m[13'd2545]=16'h000b;
m[13'd2546]=16'h0009;
m[13'd2547]=16'h110b;
m[13'd2548]=16'h0161;
m[13'd2549]=16'h0301;
m[13'd2550]=16'h0009;
m[13'd2551]=16'h9b00;
m[13'd2552]=16'h001b;
m[13'd2553]=16'h4002;
m[13'd2554]=16'h0010;
m[13'd2555]=16'h0003;
m[13'd2556]=16'h0016;
m[13'd2557]=16'h0905;
m[13'd2558]=16'h000a;
m[13'd2559]=16'h0906;
m[13'd2560]=16'h0007;
m[13'd2561]=16'h0004;
m[13'd2562]=16'h000a;
m[13'd2563]=16'h4104;
m[13'd2564]=16'h0095;
m[13'd2565]=16'h0003;
m[13'd2566]=16'h0009;
m[13'd2567]=16'h5002;
m[13'd2568]=16'h48cc;
m[13'd2569]=16'h4012;
m[13'd2570]=16'h00a0;
m[13'd2571]=16'h810b;
m[13'd2572]=16'h003b;
m[13'd2573]=16'h0808;
m[13'd2574]=16'h0009;
m[13'd2575]=16'h9307;
m[13'd2576]=16'h0072;
m[13'd2577]=16'h4801;
m[13'd2578]=16'h0007;
m[13'd2579]=16'h0000;
m[13'd2580]=16'h000e;
m[13'd2581]=16'h8104;
m[13'd2582]=16'h0060;
m[13'd2583]=16'h0003;
m[13'd2584]=16'h0009;
m[13'd2585]=16'h6002;
m[13'd2586]=16'h4af3;
m[13'd2587]=16'h4012;
m[13'd2588]=16'h00a0;
m[13'd2589]=16'h110b;
m[13'd2590]=16'h003b;
m[13'd2591]=16'h0d08;
m[13'd2592]=16'h0009;
m[13'd2593]=16'h9c07;
m[13'd2594]=16'h0090;
m[13'd2595]=16'h0301;
m[13'd2596]=16'h0009;
m[13'd2597]=16'h9b00;
m[13'd2598]=16'h0018;
m[13'd2599]=16'h4104;
m[13'd2600]=16'h0060;
m[13'd2601]=16'h0003;
m[13'd2602]=16'h0009;
m[13'd2603]=16'h7002;
m[13'd2604]=16'h4ac9;
m[13'd2605]=16'h4012;
m[13'd2606]=16'h00a0;
m[13'd2607]=16'h110b;
m[13'd2608]=16'h003b;
m[13'd2609]=16'h0a08;
m[13'd2610]=16'h0009;
m[13'd2611]=16'hcd07;
m[13'd2612]=16'h0090;
m[13'd2613]=16'h0301;
m[13'd2614]=16'h0009;
m[13'd2615]=16'h9b00;
m[13'd2616]=16'h0018;
m[13'd2617]=16'h4104;
m[13'd2618]=16'h0060;
m[13'd2619]=16'h0003;
m[13'd2620]=16'h0009;
m[13'd2621]=16'h8002;
m[13'd2622]=16'h4acc;
m[13'd2623]=16'h4012;
m[13'd2624]=16'h00a0;
m[13'd2625]=16'h100b;
m[13'd2626]=16'h003b;
m[13'd2627]=16'h0808;
m[13'd2628]=16'h0009;
m[13'd2629]=16'h9307;
m[13'd2630]=16'h0090;
m[13'd2631]=16'h0301;
m[13'd2632]=16'h0009;
m[13'd2633]=16'h9b00;
m[13'd2634]=16'h0018;
m[13'd2635]=16'h4104;
m[13'd2636]=16'h0060;
m[13'd2637]=16'h0003;
m[13'd2638]=16'h0009;
m[13'd2639]=16'h9002;
m[13'd2640]=16'h4ac9;
m[13'd2641]=16'h4012;
m[13'd2642]=16'h00a0;
m[13'd2643]=16'h100b;
m[13'd2644]=16'h003b;
m[13'd2645]=16'h0708;
m[13'd2646]=16'h0009;
m[13'd2647]=16'ha307;
m[13'd2648]=16'h0090;
m[13'd2649]=16'h0301;
m[13'd2650]=16'h0009;
m[13'd2651]=16'h9b00;
m[13'd2652]=16'h0018;
m[13'd2653]=16'h4104;
m[13'd2654]=16'h0060;
m[13'd2655]=16'h0003;
m[13'd2656]=16'h0009;
m[13'd2657]=16'ha002;
m[13'd2658]=16'h4b67;
m[13'd2659]=16'h100b;
m[13'd2660]=16'h003b;
m[13'd2661]=16'h0608;
m[13'd2662]=16'h0009;
m[13'd2663]=16'hce07;
m[13'd2664]=16'h0024;
m[13'd2665]=16'h100b;
m[13'd2666]=16'h0086;
m[13'd2667]=16'h0301;
m[13'd2668]=16'h0009;
m[13'd2669]=16'h9b00;
m[13'd2670]=16'h0018;
m[13'd2671]=16'h4104;
m[13'd2672]=16'h0025;
m[13'd2673]=16'h4004;
m[13'd2674]=16'h004e;
m[13'd2675]=16'h0003;
m[13'd2676]=16'h0009;
m[13'd2677]=16'hb002;
m[13'd2678]=16'h4b2e;
m[13'd2679]=16'h100b;
m[13'd2680]=16'h003b;
m[13'd2681]=16'h0608;
m[13'd2682]=16'h0009;
m[13'd2683]=16'h1007;
m[13'd2684]=16'h0024;
m[13'd2685]=16'h100b;
m[13'd2686]=16'h007e;
m[13'd2687]=16'h0301;
m[13'd2688]=16'h0009;
m[13'd2689]=16'h9b00;
m[13'd2690]=16'h0018;
m[13'd2691]=16'h4104;
m[13'd2692]=16'h0025;
m[13'd2693]=16'h4004;
m[13'd2694]=16'h004e;
m[13'd2695]=16'h0003;
m[13'd2696]=16'h0009;
m[13'd2697]=16'hc002;
m[13'd2698]=16'h4b45;
m[13'd2699]=16'h100b;
m[13'd2700]=16'h003a;
m[13'd2701]=16'h0508;
m[13'd2702]=16'h0009;
m[13'd2703]=16'h6707;
m[13'd2704]=16'h0024;
m[13'd2705]=16'h100b;
m[13'd2706]=16'h007e;
m[13'd2707]=16'h0301;
m[13'd2708]=16'h0009;
m[13'd2709]=16'h9b00;
m[13'd2710]=16'h0018;
m[13'd2711]=16'h4104;
m[13'd2712]=16'h0025;
m[13'd2713]=16'h4004;
m[13'd2714]=16'h004e;
m[13'd2715]=16'h0003;
m[13'd2716]=16'h0009;
m[13'd2717]=16'hd002;
m[13'd2718]=16'h4b45;
m[13'd2719]=16'h100b;
m[13'd2720]=16'h003a;
m[13'd2721]=16'h0408;
m[13'd2722]=16'h0009;
m[13'd2723]=16'hd007;
m[13'd2724]=16'h0024;
m[13'd2725]=16'h100b;
m[13'd2726]=16'h007e;
m[13'd2727]=16'h0301;
m[13'd2728]=16'h0009;
m[13'd2729]=16'h9b00;
m[13'd2730]=16'h0018;
m[13'd2731]=16'h4104;
m[13'd2732]=16'h0025;
m[13'd2733]=16'h4004;
m[13'd2734]=16'h004e;
m[13'd2735]=16'h0003;
m[13'd2736]=16'h0009;
m[13'd2737]=16'he002;
m[13'd2738]=16'h4b48;
m[13'd2739]=16'h100b;
m[13'd2740]=16'h003a;
m[13'd2741]=16'h0408;
m[13'd2742]=16'h0009;
m[13'd2743]=16'h4907;
m[13'd2744]=16'h0024;
m[13'd2745]=16'h100b;
m[13'd2746]=16'h007e;
m[13'd2747]=16'h0301;
m[13'd2748]=16'h0009;
m[13'd2749]=16'h9b00;
m[13'd2750]=16'h0018;
m[13'd2751]=16'h4104;
m[13'd2752]=16'h0025;
m[13'd2753]=16'h4004;
m[13'd2754]=16'h004e;
m[13'd2755]=16'h0003;
m[13'd2756]=16'h0009;
m[13'd2757]=16'hf002;
m[13'd2758]=16'h4b45;
m[13'd2759]=16'h100b;
m[13'd2760]=16'h003a;
m[13'd2761]=16'h0308;
m[13'd2762]=16'h0009;
m[13'd2763]=16'hd207;
m[13'd2764]=16'h0024;
m[13'd2765]=16'h100b;
m[13'd2766]=16'h007e;
m[13'd2767]=16'h0301;
m[13'd2768]=16'h0009;
m[13'd2769]=16'h9b00;
m[13'd2770]=16'h0018;
m[13'd2771]=16'h4104;
m[13'd2772]=16'h0025;
m[13'd2773]=16'h4004;
m[13'd2774]=16'h004e;
m[13'd2775]=16'h0103;
m[13'd2776]=16'h0009;
m[13'd2777]=16'h0002;
m[13'd2778]=16'h4b55;
m[13'd2779]=16'h100b;
m[13'd2780]=16'h003a;
m[13'd2781]=16'h0308;
m[13'd2782]=16'h0009;
m[13'd2783]=16'h6707;
m[13'd2784]=16'h011f;
m[13'd2785]=16'h0301;
m[13'd2786]=16'h0009;
m[13'd2787]=16'h9b00;
m[13'd2788]=16'h001b;
m[13'd2789]=16'h4002;
m[13'd2790]=16'h0010;
m[13'd2791]=16'h0003;
m[13'd2792]=16'h0016;
m[13'd2793]=16'h0905;
m[13'd2794]=16'h000a;
m[13'd2795]=16'h0906;
m[13'd2796]=16'h0007;
m[13'd2797]=16'h0004;
m[13'd2798]=16'h000a;
m[13'd2799]=16'h4104;
m[13'd2800]=16'h0095;
m[13'd2801]=16'h0003;
m[13'd2802]=16'h0009;
m[13'd2803]=16'h5002;
m[13'd2804]=16'h4a53;
m[13'd2805]=16'h000b;
m[13'd2806]=16'h003a;
m[13'd2807]=16'h0308;
m[13'd2808]=16'h0009;
m[13'd2809]=16'h6707;
m[13'd2810]=16'h0072;
m[13'd2811]=16'h4801;
m[13'd2812]=16'h0007;
m[13'd2813]=16'h0000;
m[13'd2814]=16'h000e;
m[13'd2815]=16'h8104;
m[13'd2816]=16'h0060;
m[13'd2817]=16'h0003;
m[13'd2818]=16'h0009;
m[13'd2819]=16'h6002;
m[13'd2820]=16'h4b96;
m[13'd2821]=16'h000b;
m[13'd2822]=16'h003a;
m[13'd2823]=16'h0308;
m[13'd2824]=16'h0009;
m[13'd2825]=16'h6707;
m[13'd2826]=16'h0090;
m[13'd2827]=16'h0301;
m[13'd2828]=16'h0009;
m[13'd2829]=16'h9b00;
m[13'd2830]=16'h0018;
m[13'd2831]=16'h4104;
m[13'd2832]=16'h0060;
m[13'd2833]=16'h0003;
m[13'd2834]=16'h0009;
m[13'd2835]=16'h7002;
m[13'd2836]=16'h4b6c;
m[13'd2837]=16'h000b;
m[13'd2838]=16'h003a;
m[13'd2839]=16'h0308;
m[13'd2840]=16'h0009;
m[13'd2841]=16'h6707;
m[13'd2842]=16'h0090;
m[13'd2843]=16'h0301;
m[13'd2844]=16'h0009;
m[13'd2845]=16'h9b00;
m[13'd2846]=16'h0018;
m[13'd2847]=16'h4104;
m[13'd2848]=16'h0060;
m[13'd2849]=16'h0003;
m[13'd2850]=16'h0009;
m[13'd2851]=16'h8002;
m[13'd2852]=16'h4b69;
m[13'd2853]=16'h000b;
m[13'd2854]=16'h003a;
m[13'd2855]=16'h0308;
m[13'd2856]=16'h0009;
m[13'd2857]=16'h6707;
m[13'd2858]=16'h0090;
m[13'd2859]=16'h0301;
m[13'd2860]=16'h0009;
m[13'd2861]=16'h9b00;
m[13'd2862]=16'h0018;
m[13'd2863]=16'h4104;
m[13'd2864]=16'h0060;
m[13'd2865]=16'h0003;
m[13'd2866]=16'h0009;
m[13'd2867]=16'h9002;
m[13'd2868]=16'h4b6c;
m[13'd2869]=16'h100b;
m[13'd2870]=16'h003b;
m[13'd2871]=16'h3f08;
m[13'd2872]=16'h0009;
m[13'd2873]=16'h0007;
m[13'd2874]=16'h0090;
m[13'd2875]=16'h0301;
m[13'd2876]=16'h0009;
m[13'd2877]=16'h9b00;
m[13'd2878]=16'h0018;
m[13'd2879]=16'h4104;
m[13'd2880]=16'h0060;
m[13'd2881]=16'h0003;
m[13'd2882]=16'h0009;
m[13'd2883]=16'ha002;
m[13'd2884]=16'h4bdb;
m[13'd2885]=16'h0308;
m[13'd2886]=16'h0009;
m[13'd2887]=16'h6707;
m[13'd2888]=16'h001b;
m[13'd2889]=16'h8009;
m[13'd2890]=16'h0010;
m[13'd2891]=16'h000a;
m[13'd2892]=16'h0015;
m[13'd2893]=16'h090c;
m[13'd2894]=16'h0009;
m[13'd2895]=16'h080d;
m[13'd2896]=16'h0007;
m[13'd2897]=16'h000b;
m[13'd2898]=16'h0009;
m[13'd2899]=16'h110b;
m[13'd2900]=16'h00cd;
m[13'd2901]=16'h0301;
m[13'd2902]=16'h0009;
m[13'd2903]=16'h9b00;
m[13'd2904]=16'h0018;
m[13'd2905]=16'h4104;
m[13'd2906]=16'h0025;
m[13'd2907]=16'h4004;
m[13'd2908]=16'h004e;
m[13'd2909]=16'h0003;
m[13'd2910]=16'h0009;
m[13'd2911]=16'hb002;
m[13'd2912]=16'h4a8c;
m[13'd2913]=16'h810b;
m[13'd2914]=16'h003b;
m[13'd2915]=16'h0808;
m[13'd2916]=16'h0009;
m[13'd2917]=16'h9307;
m[13'd2918]=16'h0090;
m[13'd2919]=16'h0301;
m[13'd2920]=16'h0009;
m[13'd2921]=16'h9b00;
m[13'd2922]=16'h0018;
m[13'd2923]=16'h4104;
m[13'd2924]=16'h0025;
m[13'd2925]=16'h4004;
m[13'd2926]=16'h004e;
m[13'd2927]=16'h0003;
m[13'd2928]=16'h0009;
m[13'd2929]=16'hc002;
m[13'd2930]=16'h4b57;
m[13'd2931]=16'h110b;
m[13'd2932]=16'h003b;
m[13'd2933]=16'h0d08;
m[13'd2934]=16'h0009;
m[13'd2935]=16'h9c07;
m[13'd2936]=16'h0090;
m[13'd2937]=16'h0301;
m[13'd2938]=16'h0009;
m[13'd2939]=16'h9b00;
m[13'd2940]=16'h0018;
m[13'd2941]=16'h4104;
m[13'd2942]=16'h0025;
m[13'd2943]=16'h4004;
m[13'd2944]=16'h004e;
m[13'd2945]=16'h0003;
m[13'd2946]=16'h0009;
m[13'd2947]=16'hd002;
m[13'd2948]=16'h4b57;
m[13'd2949]=16'h110b;
m[13'd2950]=16'h003b;
m[13'd2951]=16'h0a08;
m[13'd2952]=16'h0009;
m[13'd2953]=16'hcd07;
m[13'd2954]=16'h0090;
m[13'd2955]=16'h0301;
m[13'd2956]=16'h0009;
m[13'd2957]=16'h9b00;
m[13'd2958]=16'h0018;
m[13'd2959]=16'h4104;
m[13'd2960]=16'h0025;
m[13'd2961]=16'h4004;
m[13'd2962]=16'h004e;
m[13'd2963]=16'h0003;
m[13'd2964]=16'h0009;
m[13'd2965]=16'he002;
m[13'd2966]=16'h4b57;
m[13'd2967]=16'h100b;
m[13'd2968]=16'h003b;
m[13'd2969]=16'h0808;
m[13'd2970]=16'h0009;
m[13'd2971]=16'h9307;
m[13'd2972]=16'h0090;
m[13'd2973]=16'h0301;
m[13'd2974]=16'h0009;
m[13'd2975]=16'h9b00;
m[13'd2976]=16'h0018;
m[13'd2977]=16'h4104;
m[13'd2978]=16'h0025;
m[13'd2979]=16'h4004;
m[13'd2980]=16'h004e;
m[13'd2981]=16'h0003;
m[13'd2982]=16'h0009;
m[13'd2983]=16'hf002;
m[13'd2984]=16'h4b57;
m[13'd2985]=16'h100b;
m[13'd2986]=16'h003b;
m[13'd2987]=16'h0708;
m[13'd2988]=16'h0009;
m[13'd2989]=16'ha307;
m[13'd2990]=16'h0090;
m[13'd2991]=16'h0301;
m[13'd2992]=16'h0009;
m[13'd2993]=16'h9b00;
m[13'd2994]=16'h0018;
m[13'd2995]=16'h4104;
m[13'd2996]=16'h0025;
m[13'd2997]=16'h4004;
m[13'd2998]=16'h004e;
m[13'd2999]=16'h0103;
m[13'd3000]=16'h0009;
m[13'd3001]=16'h0002;
m[13'd3002]=16'h4b67;
m[13'd3003]=16'h100b;
m[13'd3004]=16'h003b;
m[13'd3005]=16'h0608;
m[13'd3006]=16'h0009;
m[13'd3007]=16'hce07;
m[13'd3008]=16'h0024;
m[13'd3009]=16'h100b;
m[13'd3010]=16'h011a;
m[13'd3011]=16'h0301;
m[13'd3012]=16'h0009;
m[13'd3013]=16'h9b00;
m[13'd3014]=16'h001b;
m[13'd3015]=16'h4002;
m[13'd3016]=16'h0010;
m[13'd3017]=16'h0003;
m[13'd3018]=16'h0016;
m[13'd3019]=16'h0905;
m[13'd3020]=16'h000a;
m[13'd3021]=16'h0906;
m[13'd3022]=16'h0007;
m[13'd3023]=16'h0004;
m[13'd3024]=16'h000a;
m[13'd3025]=16'h4104;
m[13'd3026]=16'h008d;
m[13'd3027]=16'h0003;
m[13'd3028]=16'h0009;
m[13'd3029]=16'h5002;
m[13'd3030]=16'h4a3b;
m[13'd3031]=16'h100b;
m[13'd3032]=16'h003b;
m[13'd3033]=16'h0608;
m[13'd3034]=16'h0009;
m[13'd3035]=16'h1007;
m[13'd3036]=16'h0024;
m[13'd3037]=16'h100b;
m[13'd3038]=16'h0060;
m[13'd3039]=16'h4801;
m[13'd3040]=16'h0007;
m[13'd3041]=16'h0000;
m[13'd3042]=16'h000e;
m[13'd3043]=16'h8104;
m[13'd3044]=16'h0058;
m[13'd3045]=16'h0003;
m[13'd3046]=16'h0009;
m[13'd3047]=16'h6002;
m[13'd3048]=16'h4b8a;
m[13'd3049]=16'h100b;
m[13'd3050]=16'h003a;
m[13'd3051]=16'h0508;
m[13'd3052]=16'h0009;
m[13'd3053]=16'h6707;
m[13'd3054]=16'h0024;
m[13'd3055]=16'h100b;
m[13'd3056]=16'h007e;
m[13'd3057]=16'h0301;
m[13'd3058]=16'h0009;
m[13'd3059]=16'h9b00;
m[13'd3060]=16'h0018;
m[13'd3061]=16'h4104;
m[13'd3062]=16'h0058;
m[13'd3063]=16'h0003;
m[13'd3064]=16'h0009;
m[13'd3065]=16'h7002;
m[13'd3066]=16'h4b60;
m[13'd3067]=16'h100b;
m[13'd3068]=16'h003a;
m[13'd3069]=16'h0408;
m[13'd3070]=16'h0009;
m[13'd3071]=16'hd007;
m[13'd3072]=16'h0024;
m[13'd3073]=16'h100b;
m[13'd3074]=16'h007e;
m[13'd3075]=16'h0301;
m[13'd3076]=16'h0009;
m[13'd3077]=16'h9b00;
m[13'd3078]=16'h0018;
m[13'd3079]=16'h4104;
m[13'd3080]=16'h0058;
m[13'd3081]=16'h0003;
m[13'd3082]=16'h0009;
m[13'd3083]=16'h8002;
m[13'd3084]=16'h4b60;
m[13'd3085]=16'h100b;
m[13'd3086]=16'h003a;
m[13'd3087]=16'h0408;
m[13'd3088]=16'h0009;
m[13'd3089]=16'h4907;
m[13'd3090]=16'h0024;
m[13'd3091]=16'h100b;
m[13'd3092]=16'h007e;
m[13'd3093]=16'h0301;
m[13'd3094]=16'h0009;
m[13'd3095]=16'h9b00;
m[13'd3096]=16'h0018;
m[13'd3097]=16'h4104;
m[13'd3098]=16'h0058;
m[13'd3099]=16'h0003;
m[13'd3100]=16'h0009;
m[13'd3101]=16'h9002;
m[13'd3102]=16'h4b63;
m[13'd3103]=16'h100b;
m[13'd3104]=16'h003a;
m[13'd3105]=16'h0308;
m[13'd3106]=16'h0009;
m[13'd3107]=16'hd207;
m[13'd3108]=16'h0024;
m[13'd3109]=16'h100b;
m[13'd3110]=16'h007e;
m[13'd3111]=16'h0301;
m[13'd3112]=16'h0009;
m[13'd3113]=16'h9b00;
m[13'd3114]=16'h0018;
m[13'd3115]=16'h4104;
m[13'd3116]=16'h0058;
m[13'd3117]=16'h0003;
m[13'd3118]=16'h0009;
m[13'd3119]=16'ha002;
m[13'd3120]=16'h4b70;
m[13'd3121]=16'h100b;
m[13'd3122]=16'h003a;
m[13'd3123]=16'h0308;
m[13'd3124]=16'h0009;
m[13'd3125]=16'h6707;
m[13'd3126]=16'h011f;
m[13'd3127]=16'h0401;
m[13'd3128]=16'h0009;
m[13'd3129]=16'h4900;
m[13'd3130]=16'h001b;
m[13'd3131]=16'h4002;
m[13'd3132]=16'h0010;
m[13'd3133]=16'h0003;
m[13'd3134]=16'h0016;
m[13'd3135]=16'h0905;
m[13'd3136]=16'h000a;
m[13'd3137]=16'h0906;
m[13'd3138]=16'h0007;
m[13'd3139]=16'h0004;
m[13'd3140]=16'h000a;
m[13'd3141]=16'h4104;
m[13'd3142]=16'h008d;
m[13'd3143]=16'h0003;
m[13'd3144]=16'h0009;
m[13'd3145]=16'h5002;
m[13'd3146]=16'h4a5c;
m[13'd3147]=16'h000b;
m[13'd3148]=16'h003a;
m[13'd3149]=16'h0308;
m[13'd3150]=16'h0009;
m[13'd3151]=16'h6707;
m[13'd3152]=16'h0072;
m[13'd3153]=16'h4801;
m[13'd3154]=16'h0007;
m[13'd3155]=16'h0000;
m[13'd3156]=16'h000e;
m[13'd3157]=16'h8104;
m[13'd3158]=16'h0058;
m[13'd3159]=16'h0003;
m[13'd3160]=16'h0009;
m[13'd3161]=16'h6002;
m[13'd3162]=16'h4b9c;
m[13'd3163]=16'h000b;
m[13'd3164]=16'h003a;
m[13'd3165]=16'h0308;
m[13'd3166]=16'h0009;
m[13'd3167]=16'h6707;
m[13'd3168]=16'h0090;
m[13'd3169]=16'h0401;
m[13'd3170]=16'h0009;
m[13'd3171]=16'h4900;
m[13'd3172]=16'h0018;
m[13'd3173]=16'h4104;
m[13'd3174]=16'h0058;
m[13'd3175]=16'h0003;
m[13'd3176]=16'h0009;
m[13'd3177]=16'h7002;
m[13'd3178]=16'h4b72;
m[13'd3179]=16'h000b;
m[13'd3180]=16'h003a;
m[13'd3181]=16'h0308;
m[13'd3182]=16'h0009;
m[13'd3183]=16'h6707;
m[13'd3184]=16'h0090;
m[13'd3185]=16'h0401;
m[13'd3186]=16'h0009;
m[13'd3187]=16'h4900;
m[13'd3188]=16'h0018;
m[13'd3189]=16'h4104;
m[13'd3190]=16'h0058;
m[13'd3191]=16'h0003;
m[13'd3192]=16'h0009;
m[13'd3193]=16'h8002;
m[13'd3194]=16'h4b75;
m[13'd3195]=16'h000b;
m[13'd3196]=16'h003a;
m[13'd3197]=16'h0308;
m[13'd3198]=16'h0009;
m[13'd3199]=16'h6707;
m[13'd3200]=16'h0090;
m[13'd3201]=16'h0401;
m[13'd3202]=16'h0009;
m[13'd3203]=16'h4900;
m[13'd3204]=16'h0018;
m[13'd3205]=16'h4104;
m[13'd3206]=16'h0058;
m[13'd3207]=16'h0003;
m[13'd3208]=16'h0009;
m[13'd3209]=16'h9002;
m[13'd3210]=16'h4b72;
m[13'd3211]=16'h100b;
m[13'd3212]=16'h003b;
m[13'd3213]=16'h3f08;
m[13'd3214]=16'h0009;
m[13'd3215]=16'h0007;
m[13'd3216]=16'h0090;
m[13'd3217]=16'h0401;
m[13'd3218]=16'h0009;
m[13'd3219]=16'h4900;
m[13'd3220]=16'h0018;
m[13'd3221]=16'h4104;
m[13'd3222]=16'h0058;
m[13'd3223]=16'h0003;
m[13'd3224]=16'h0009;
m[13'd3225]=16'ha002;
m[13'd3226]=16'h4be4;
m[13'd3227]=16'h0308;
m[13'd3228]=16'h0009;
m[13'd3229]=16'h6707;
m[13'd3230]=16'h001b;
m[13'd3231]=16'h8009;
m[13'd3232]=16'h0010;
m[13'd3233]=16'h000a;
m[13'd3234]=16'h0015;
m[13'd3235]=16'h090c;
m[13'd3236]=16'h0009;
m[13'd3237]=16'h080d;
m[13'd3238]=16'h0007;
m[13'd3239]=16'h000b;
m[13'd3240]=16'h0009;
m[13'd3241]=16'h110b;
m[13'd3242]=16'h0161;
m[13'd3243]=16'h0301;
m[13'd3244]=16'h0009;
m[13'd3245]=16'h9b00;
m[13'd3246]=16'h001b;
m[13'd3247]=16'h4002;
m[13'd3248]=16'h0010;
m[13'd3249]=16'h0003;
m[13'd3250]=16'h0016;
m[13'd3251]=16'h0905;
m[13'd3252]=16'h000a;
m[13'd3253]=16'h0906;
m[13'd3254]=16'h0007;
m[13'd3255]=16'h0004;
m[13'd3256]=16'h000a;
m[13'd3257]=16'h4104;
m[13'd3258]=16'h0095;
m[13'd3259]=16'h0003;
m[13'd3260]=16'h0009;
m[13'd3261]=16'h5002;
m[13'd3262]=16'h4990;
m[13'd3263]=16'h810b;
m[13'd3264]=16'h003b;
m[13'd3265]=16'h0808;
m[13'd3266]=16'h0009;
m[13'd3267]=16'h9307;
m[13'd3268]=16'h0072;
m[13'd3269]=16'h4801;
m[13'd3270]=16'h0007;
m[13'd3271]=16'h0000;
m[13'd3272]=16'h000e;
m[13'd3273]=16'h8104;
m[13'd3274]=16'h0060;
m[13'd3275]=16'h0003;
m[13'd3276]=16'h0009;
m[13'd3277]=16'h6002;
m[13'd3278]=16'h4b93;
m[13'd3279]=16'h110b;
m[13'd3280]=16'h003b;
m[13'd3281]=16'h0d08;
m[13'd3282]=16'h0009;
m[13'd3283]=16'h9c07;
m[13'd3284]=16'h0090;
m[13'd3285]=16'h0301;
m[13'd3286]=16'h0009;
m[13'd3287]=16'h9b00;
m[13'd3288]=16'h0018;
m[13'd3289]=16'h4104;
m[13'd3290]=16'h0060;
m[13'd3291]=16'h0003;
m[13'd3292]=16'h0009;
m[13'd3293]=16'h7002;
m[13'd3294]=16'h4b6c;
m[13'd3295]=16'h110b;
m[13'd3296]=16'h003b;
m[13'd3297]=16'h0a08;
m[13'd3298]=16'h0009;
m[13'd3299]=16'hcd07;
m[13'd3300]=16'h0090;
m[13'd3301]=16'h0301;
m[13'd3302]=16'h0009;
m[13'd3303]=16'h9b00;
m[13'd3304]=16'h0018;
m[13'd3305]=16'h4104;
m[13'd3306]=16'h0060;
m[13'd3307]=16'h0003;
m[13'd3308]=16'h0009;
m[13'd3309]=16'h8002;
m[13'd3310]=16'h4b69;
m[13'd3311]=16'h100b;
m[13'd3312]=16'h003b;
m[13'd3313]=16'h0808;
m[13'd3314]=16'h0009;
m[13'd3315]=16'h9307;
m[13'd3316]=16'h0090;
m[13'd3317]=16'h0301;
m[13'd3318]=16'h0009;
m[13'd3319]=16'h9b00;
m[13'd3320]=16'h0018;
m[13'd3321]=16'h4104;
m[13'd3322]=16'h0060;
m[13'd3323]=16'h0003;
m[13'd3324]=16'h0009;
m[13'd3325]=16'h9002;
m[13'd3326]=16'h4b69;
m[13'd3327]=16'h100b;
m[13'd3328]=16'h003b;
m[13'd3329]=16'h0708;
m[13'd3330]=16'h0009;
m[13'd3331]=16'ha307;
m[13'd3332]=16'h0090;
m[13'd3333]=16'h0301;
m[13'd3334]=16'h0009;
m[13'd3335]=16'h9b00;
m[13'd3336]=16'h0018;
m[13'd3337]=16'h4104;
m[13'd3338]=16'h0060;
m[13'd3339]=16'h0003;
m[13'd3340]=16'h0009;
m[13'd3341]=16'ha002;
m[13'd3342]=16'h4b7c;
m[13'd3343]=16'h100b;
m[13'd3344]=16'h003b;
m[13'd3345]=16'h0608;
m[13'd3346]=16'h0009;
m[13'd3347]=16'hce07;
m[13'd3348]=16'h0024;
m[13'd3349]=16'h100b;
m[13'd3350]=16'h0086;
m[13'd3351]=16'h0301;
m[13'd3352]=16'h0009;
m[13'd3353]=16'h9b00;
m[13'd3354]=16'h0018;
m[13'd3355]=16'h4104;
m[13'd3356]=16'h0025;
m[13'd3357]=16'h4004;
m[13'd3358]=16'h004e;
m[13'd3359]=16'h0003;
m[13'd3360]=16'h0009;
m[13'd3361]=16'hb002;
m[13'd3362]=16'h4b2b;
m[13'd3363]=16'h100b;
m[13'd3364]=16'h003b;
m[13'd3365]=16'h0608;
m[13'd3366]=16'h0009;
m[13'd3367]=16'h1007;
m[13'd3368]=16'h0024;
m[13'd3369]=16'h100b;
m[13'd3370]=16'h007e;
m[13'd3371]=16'h0301;
m[13'd3372]=16'h0009;
m[13'd3373]=16'h9b00;
m[13'd3374]=16'h0018;
m[13'd3375]=16'h4104;
m[13'd3376]=16'h0025;
m[13'd3377]=16'h4004;
m[13'd3378]=16'h004e;
m[13'd3379]=16'h0003;
m[13'd3380]=16'h0009;
m[13'd3381]=16'hc002;
m[13'd3382]=16'h4b45;
m[13'd3383]=16'h100b;
m[13'd3384]=16'h003a;
m[13'd3385]=16'h0508;
m[13'd3386]=16'h0009;
m[13'd3387]=16'h6707;
m[13'd3388]=16'h0024;
m[13'd3389]=16'h100b;
m[13'd3390]=16'h007e;
m[13'd3391]=16'h0301;
m[13'd3392]=16'h0009;
m[13'd3393]=16'h9b00;
m[13'd3394]=16'h0018;
m[13'd3395]=16'h4104;
m[13'd3396]=16'h0025;
m[13'd3397]=16'h4004;
m[13'd3398]=16'h004e;
m[13'd3399]=16'h0003;
m[13'd3400]=16'h0009;
m[13'd3401]=16'hd002;
m[13'd3402]=16'h4b48;
m[13'd3403]=16'h100b;
m[13'd3404]=16'h003a;
m[13'd3405]=16'h0408;
m[13'd3406]=16'h0009;
m[13'd3407]=16'hd007;
m[13'd3408]=16'h0024;
m[13'd3409]=16'h100b;
m[13'd3410]=16'h007e;
m[13'd3411]=16'h0301;
m[13'd3412]=16'h0009;
m[13'd3413]=16'h9b00;
m[13'd3414]=16'h0018;
m[13'd3415]=16'h4104;
m[13'd3416]=16'h0025;
m[13'd3417]=16'h4004;
m[13'd3418]=16'h004e;
m[13'd3419]=16'h0003;
m[13'd3420]=16'h0009;
m[13'd3421]=16'he002;
m[13'd3422]=16'h4b45;
m[13'd3423]=16'h100b;
m[13'd3424]=16'h003a;
m[13'd3425]=16'h0408;
m[13'd3426]=16'h0009;
m[13'd3427]=16'h4907;
m[13'd3428]=16'h0024;
m[13'd3429]=16'h100b;
m[13'd3430]=16'h007e;
m[13'd3431]=16'h0301;
m[13'd3432]=16'h0009;
m[13'd3433]=16'h9b00;
m[13'd3434]=16'h0018;
m[13'd3435]=16'h4104;
m[13'd3436]=16'h0025;
m[13'd3437]=16'h4004;
m[13'd3438]=16'h004e;
m[13'd3439]=16'h0003;
m[13'd3440]=16'h0009;
m[13'd3441]=16'hf002;
m[13'd3442]=16'h4b45;
m[13'd3443]=16'h100b;
m[13'd3444]=16'h003a;
m[13'd3445]=16'h0308;
m[13'd3446]=16'h0009;
m[13'd3447]=16'hd207;
m[13'd3448]=16'h0024;
m[13'd3449]=16'h100b;
m[13'd3450]=16'h007e;
m[13'd3451]=16'h0301;
m[13'd3452]=16'h0009;
m[13'd3453]=16'h9b00;
m[13'd3454]=16'h0018;
m[13'd3455]=16'h4104;
m[13'd3456]=16'h0025;
m[13'd3457]=16'h4004;
m[13'd3458]=16'h004e;
m[13'd3459]=16'h0103;
m[13'd3460]=16'h0009;
m[13'd3461]=16'h0002;
m[13'd3462]=16'h4b58;
m[13'd3463]=16'h100b;
m[13'd3464]=16'h003a;
m[13'd3465]=16'h0308;
m[13'd3466]=16'h0009;
m[13'd3467]=16'h6707;
m[13'd3468]=16'h012c;
m[13'd3469]=16'h0401;
m[13'd3470]=16'h0009;
m[13'd3471]=16'hd000;
m[13'd3472]=16'h001b;
m[13'd3473]=16'h4002;
m[13'd3474]=16'h0010;
m[13'd3475]=16'h0003;
m[13'd3476]=16'h0016;
m[13'd3477]=16'h0905;
m[13'd3478]=16'h000a;
m[13'd3479]=16'h0906;
m[13'd3480]=16'h0007;
m[13'd3481]=16'h0004;
m[13'd3482]=16'h000a;
m[13'd3483]=16'h4104;
m[13'd3484]=16'h008d;
m[13'd3485]=16'h0003;
m[13'd3486]=16'h0009;
m[13'd3487]=16'h5002;
m[13'd3488]=16'h4a4d;
m[13'd3489]=16'h000b;
m[13'd3490]=16'h003a;
m[13'd3491]=16'h0308;
m[13'd3492]=16'h0009;
m[13'd3493]=16'h6707;
m[13'd3494]=16'h0072;
m[13'd3495]=16'h4801;
m[13'd3496]=16'h0007;
m[13'd3497]=16'h0000;
m[13'd3498]=16'h000e;
m[13'd3499]=16'h8104;
m[13'd3500]=16'h0058;
m[13'd3501]=16'h0003;
m[13'd3502]=16'h0009;
m[13'd3503]=16'h6002;
m[13'd3504]=16'h4b9c;
m[13'd3505]=16'h000b;
m[13'd3506]=16'h003a;
m[13'd3507]=16'h0308;
m[13'd3508]=16'h0009;
m[13'd3509]=16'h6707;
m[13'd3510]=16'h0090;
m[13'd3511]=16'h0401;
m[13'd3512]=16'h0009;
m[13'd3513]=16'hd000;
m[13'd3514]=16'h0018;
m[13'd3515]=16'h4104;
m[13'd3516]=16'h0058;
m[13'd3517]=16'h0003;
m[13'd3518]=16'h0009;
m[13'd3519]=16'h7002;
m[13'd3520]=16'h4b75;
m[13'd3521]=16'h000b;
m[13'd3522]=16'h003a;
m[13'd3523]=16'h0308;
m[13'd3524]=16'h0009;
m[13'd3525]=16'h6707;
m[13'd3526]=16'h0090;
m[13'd3527]=16'h0401;
m[13'd3528]=16'h0009;
m[13'd3529]=16'hd000;
m[13'd3530]=16'h0018;
m[13'd3531]=16'h4104;
m[13'd3532]=16'h0058;
m[13'd3533]=16'h0003;
m[13'd3534]=16'h0009;
m[13'd3535]=16'h8002;
m[13'd3536]=16'h4b72;
m[13'd3537]=16'h000b;
m[13'd3538]=16'h003a;
m[13'd3539]=16'h0308;
m[13'd3540]=16'h0009;
m[13'd3541]=16'h6707;
m[13'd3542]=16'h0090;
m[13'd3543]=16'h0401;
m[13'd3544]=16'h0009;
m[13'd3545]=16'hd000;
m[13'd3546]=16'h0018;
m[13'd3547]=16'h4104;
m[13'd3548]=16'h0058;
m[13'd3549]=16'h0003;
m[13'd3550]=16'h0009;
m[13'd3551]=16'h9002;
m[13'd3552]=16'h4b72;
m[13'd3553]=16'h100b;
m[13'd3554]=16'h003b;
m[13'd3555]=16'h3f08;
m[13'd3556]=16'h0009;
m[13'd3557]=16'h0007;
m[13'd3558]=16'h0090;
m[13'd3559]=16'h0401;
m[13'd3560]=16'h0009;
m[13'd3561]=16'hd000;
m[13'd3562]=16'h0018;
m[13'd3563]=16'h4104;
m[13'd3564]=16'h0058;
m[13'd3565]=16'h0003;
m[13'd3566]=16'h0009;
m[13'd3567]=16'ha002;
m[13'd3568]=16'h4bf1;
m[13'd3569]=16'h0308;
m[13'd3570]=16'h0009;
m[13'd3571]=16'h6707;
m[13'd3572]=16'h001b;
m[13'd3573]=16'h8009;
m[13'd3574]=16'h0010;
m[13'd3575]=16'h000a;
m[13'd3576]=16'h0015;
m[13'd3577]=16'h090c;
m[13'd3578]=16'h0009;
m[13'd3579]=16'h080d;
m[13'd3580]=16'h0007;
m[13'd3581]=16'h000b;
m[13'd3582]=16'h0009;
m[13'd3583]=16'h110b;
m[13'd3584]=16'h0154;
m[13'd3585]=16'h0501;
m[13'd3586]=16'h0009;
m[13'd3587]=16'h1900;
m[13'd3588]=16'h001b;
m[13'd3589]=16'h4002;
m[13'd3590]=16'h0010;
m[13'd3591]=16'h0003;
m[13'd3592]=16'h0016;
m[13'd3593]=16'h0905;
m[13'd3594]=16'h000a;
m[13'd3595]=16'h0906;
m[13'd3596]=16'h0007;
m[13'd3597]=16'h0004;
m[13'd3598]=16'h000a;
m[13'd3599]=16'h4104;
m[13'd3600]=16'h008d;
m[13'd3601]=16'h0003;
m[13'd3602]=16'h0009;
m[13'd3603]=16'h5002;
m[13'd3604]=16'h4999;
m[13'd3605]=16'h810b;
m[13'd3606]=16'h003b;
m[13'd3607]=16'h0808;
m[13'd3608]=16'h0009;
m[13'd3609]=16'h9307;
m[13'd3610]=16'h0072;
m[13'd3611]=16'h4801;
m[13'd3612]=16'h0007;
m[13'd3613]=16'h0000;
m[13'd3614]=16'h000e;
m[13'd3615]=16'h8104;
m[13'd3616]=16'h0058;
m[13'd3617]=16'h0003;
m[13'd3618]=16'h0009;
m[13'd3619]=16'h6002;
m[13'd3620]=16'h4b9c;
m[13'd3621]=16'h110b;
m[13'd3622]=16'h003b;
m[13'd3623]=16'h0d08;
m[13'd3624]=16'h0009;
m[13'd3625]=16'h9c07;
m[13'd3626]=16'h0090;
m[13'd3627]=16'h0501;
m[13'd3628]=16'h0009;
m[13'd3629]=16'h1900;
m[13'd3630]=16'h0018;
m[13'd3631]=16'h4104;
m[13'd3632]=16'h0058;
m[13'd3633]=16'h0003;
m[13'd3634]=16'h0009;
m[13'd3635]=16'h7002;
m[13'd3636]=16'h4b72;
m[13'd3637]=16'h110b;
m[13'd3638]=16'h003b;
m[13'd3639]=16'h0a08;
m[13'd3640]=16'h0009;
m[13'd3641]=16'hcd07;
m[13'd3642]=16'h0090;
m[13'd3643]=16'h0501;
m[13'd3644]=16'h0009;
m[13'd3645]=16'h1900;
m[13'd3646]=16'h0018;
m[13'd3647]=16'h4104;
m[13'd3648]=16'h0058;
m[13'd3649]=16'h0003;
m[13'd3650]=16'h0009;
m[13'd3651]=16'h8002;
m[13'd3652]=16'h4b72;
m[13'd3653]=16'h100b;
m[13'd3654]=16'h003b;
m[13'd3655]=16'h0808;
m[13'd3656]=16'h0009;
m[13'd3657]=16'h9307;
m[13'd3658]=16'h0090;
m[13'd3659]=16'h0501;
m[13'd3660]=16'h0009;
m[13'd3661]=16'h1900;
m[13'd3662]=16'h0018;
m[13'd3663]=16'h4104;
m[13'd3664]=16'h0058;
m[13'd3665]=16'h0003;
m[13'd3666]=16'h0009;
m[13'd3667]=16'h9002;
m[13'd3668]=16'h4b72;
m[13'd3669]=16'h100b;
m[13'd3670]=16'h003b;
m[13'd3671]=16'h0708;
m[13'd3672]=16'h0009;
m[13'd3673]=16'ha307;
m[13'd3674]=16'h0090;
m[13'd3675]=16'h0501;
m[13'd3676]=16'h0009;
m[13'd3677]=16'h1900;
m[13'd3678]=16'h0018;
m[13'd3679]=16'h4104;
m[13'd3680]=16'h0058;
m[13'd3681]=16'h0003;
m[13'd3682]=16'h0009;
m[13'd3683]=16'ha002;
m[13'd3684]=16'h4b82;
m[13'd3685]=16'h100b;
m[13'd3686]=16'h003b;
m[13'd3687]=16'h0608;
m[13'd3688]=16'h0009;
m[13'd3689]=16'hce07;
m[13'd3690]=16'h0024;
m[13'd3691]=16'h100b;
m[13'd3692]=16'h010d;
m[13'd3693]=16'h0501;
m[13'd3694]=16'h0009;
m[13'd3695]=16'h6700;
m[13'd3696]=16'h001b;
m[13'd3697]=16'h4002;
m[13'd3698]=16'h0010;
m[13'd3699]=16'h0003;
m[13'd3700]=16'h0016;
m[13'd3701]=16'h0905;
m[13'd3702]=16'h000a;
m[13'd3703]=16'h0906;
m[13'd3704]=16'h0007;
m[13'd3705]=16'h0004;
m[13'd3706]=16'h000a;
m[13'd3707]=16'h4104;
m[13'd3708]=16'h008d;
m[13'd3709]=16'h0003;
m[13'd3710]=16'h0009;
m[13'd3711]=16'h5002;
m[13'd3712]=16'h4a47;
m[13'd3713]=16'h100b;
m[13'd3714]=16'h003b;
m[13'd3715]=16'h0608;
m[13'd3716]=16'h0009;
m[13'd3717]=16'h1007;
m[13'd3718]=16'h0024;
m[13'd3719]=16'h100b;
m[13'd3720]=16'h0060;
m[13'd3721]=16'h4801;
m[13'd3722]=16'h0007;
m[13'd3723]=16'h0000;
m[13'd3724]=16'h000e;
m[13'd3725]=16'h8104;
m[13'd3726]=16'h0058;
m[13'd3727]=16'h0003;
m[13'd3728]=16'h0009;
m[13'd3729]=16'h6002;
m[13'd3730]=16'h4b8a;
m[13'd3731]=16'h100b;
m[13'd3732]=16'h003a;
m[13'd3733]=16'h0508;
m[13'd3734]=16'h0009;
m[13'd3735]=16'h6707;
m[13'd3736]=16'h0024;
m[13'd3737]=16'h100b;
m[13'd3738]=16'h007e;
m[13'd3739]=16'h0501;
m[13'd3740]=16'h0009;
m[13'd3741]=16'h6700;
m[13'd3742]=16'h0018;
m[13'd3743]=16'h4104;
m[13'd3744]=16'h0058;
m[13'd3745]=16'h0003;
m[13'd3746]=16'h0009;
m[13'd3747]=16'h7002;
m[13'd3748]=16'h4b63;
m[13'd3749]=16'h100b;
m[13'd3750]=16'h003a;
m[13'd3751]=16'h0408;
m[13'd3752]=16'h0009;
m[13'd3753]=16'hd007;
m[13'd3754]=16'h0024;
m[13'd3755]=16'h100b;
m[13'd3756]=16'h007e;
m[13'd3757]=16'h0501;
m[13'd3758]=16'h0009;
m[13'd3759]=16'h6700;
m[13'd3760]=16'h0018;
m[13'd3761]=16'h4104;
m[13'd3762]=16'h0058;
m[13'd3763]=16'h0003;
m[13'd3764]=16'h0009;
m[13'd3765]=16'h8002;
m[13'd3766]=16'h4b60;
m[13'd3767]=16'h100b;
m[13'd3768]=16'h003a;
m[13'd3769]=16'h0408;
m[13'd3770]=16'h0009;
m[13'd3771]=16'h4907;
m[13'd3772]=16'h0024;
m[13'd3773]=16'h100b;
m[13'd3774]=16'h007e;
m[13'd3775]=16'h0501;
m[13'd3776]=16'h0009;
m[13'd3777]=16'h6700;
m[13'd3778]=16'h0018;
m[13'd3779]=16'h4104;
m[13'd3780]=16'h0058;
m[13'd3781]=16'h0003;
m[13'd3782]=16'h0009;
m[13'd3783]=16'h9002;
m[13'd3784]=16'h4b60;
m[13'd3785]=16'h100b;
m[13'd3786]=16'h003a;
m[13'd3787]=16'h0308;
m[13'd3788]=16'h0009;
m[13'd3789]=16'hd207;
m[13'd3790]=16'h0024;
m[13'd3791]=16'h100b;
m[13'd3792]=16'h007e;
m[13'd3793]=16'h0501;
m[13'd3794]=16'h0009;
m[13'd3795]=16'h6700;
m[13'd3796]=16'h0018;
m[13'd3797]=16'h4104;
m[13'd3798]=16'h0058;
m[13'd3799]=16'h0003;
m[13'd3800]=16'h0009;
m[13'd3801]=16'ha002;
m[13'd3802]=16'h4be2;
m[13'd3803]=16'h0308;
m[13'd3804]=16'h0009;
m[13'd3805]=16'h6707;
m[13'd3806]=16'h001b;
m[13'd3807]=16'h8009;
m[13'd3808]=16'h0010;
m[13'd3809]=16'h000a;
m[13'd3810]=16'h0015;
m[13'd3811]=16'h090c;
m[13'd3812]=16'h0009;
m[13'd3813]=16'h080d;
m[13'd3814]=16'h0007;
m[13'd3815]=16'h000b;
m[13'd3816]=16'h0009;
m[13'd3817]=16'h110b;
m[13'd3818]=16'h015a;
m[13'd3819]=16'h0601;
m[13'd3820]=16'h0009;
m[13'd3821]=16'h6c00;
m[13'd3822]=16'h001b;
m[13'd3823]=16'h4002;
m[13'd3824]=16'h0010;
m[13'd3825]=16'h0003;
m[13'd3826]=16'h0016;
m[13'd3827]=16'h0905;
m[13'd3828]=16'h000a;
m[13'd3829]=16'h0906;
m[13'd3830]=16'h0007;
m[13'd3831]=16'h0004;
m[13'd3832]=16'h000a;
m[13'd3833]=16'h4104;
m[13'd3834]=16'h0095;
m[13'd3835]=16'h0003;
m[13'd3836]=16'h0009;
m[13'd3837]=16'h5002;
m[13'd3838]=16'h498a;
m[13'd3839]=16'h810b;
m[13'd3840]=16'h003b;
m[13'd3841]=16'h0808;
m[13'd3842]=16'h0009;
m[13'd3843]=16'h9307;
m[13'd3844]=16'h006a;
m[13'd3845]=16'h4801;
m[13'd3846]=16'h0007;
m[13'd3847]=16'h0000;
m[13'd3848]=16'h000e;
m[13'd3849]=16'h8104;
m[13'd3850]=16'h0060;
m[13'd3851]=16'h0003;
m[13'd3852]=16'h0009;
m[13'd3853]=16'h6002;
m[13'd3854]=16'h4b9c;
m[13'd3855]=16'h110b;
m[13'd3856]=16'h003b;
m[13'd3857]=16'h0d08;
m[13'd3858]=16'h0009;
m[13'd3859]=16'h9c07;
m[13'd3860]=16'h0089;
m[13'd3861]=16'h0601;
m[13'd3862]=16'h0009;
m[13'd3863]=16'h6c00;
m[13'd3864]=16'h0018;
m[13'd3865]=16'h4104;
m[13'd3866]=16'h0060;
m[13'd3867]=16'h0003;
m[13'd3868]=16'h0009;
m[13'd3869]=16'h7002;
m[13'd3870]=16'h4b6f;
m[13'd3871]=16'h110b;
m[13'd3872]=16'h003b;
m[13'd3873]=16'h0a08;
m[13'd3874]=16'h0009;
m[13'd3875]=16'hcd07;
m[13'd3876]=16'h0089;
m[13'd3877]=16'h0601;
m[13'd3878]=16'h0009;
m[13'd3879]=16'h6c00;
m[13'd3880]=16'h0018;
m[13'd3881]=16'h4104;
m[13'd3882]=16'h0060;
m[13'd3883]=16'h0003;
m[13'd3884]=16'h0009;
m[13'd3885]=16'h8002;
m[13'd3886]=16'h4b72;
m[13'd3887]=16'h100b;
m[13'd3888]=16'h003b;
m[13'd3889]=16'h0808;
m[13'd3890]=16'h0009;
m[13'd3891]=16'h9307;
m[13'd3892]=16'h0089;
m[13'd3893]=16'h0601;
m[13'd3894]=16'h0009;
m[13'd3895]=16'h6c00;
m[13'd3896]=16'h0018;
m[13'd3897]=16'h4104;
m[13'd3898]=16'h0060;
m[13'd3899]=16'h0003;
m[13'd3900]=16'h0009;
m[13'd3901]=16'h9002;
m[13'd3902]=16'h4b72;
m[13'd3903]=16'h100b;
m[13'd3904]=16'h003b;
m[13'd3905]=16'h0708;
m[13'd3906]=16'h0009;
m[13'd3907]=16'ha307;
m[13'd3908]=16'h0089;
m[13'd3909]=16'h0601;
m[13'd3910]=16'h0009;
m[13'd3911]=16'h6c00;
m[13'd3912]=16'h0018;
m[13'd3913]=16'h4104;
m[13'd3914]=16'h0060;
m[13'd3915]=16'h0003;
m[13'd3916]=16'h0009;
m[13'd3917]=16'ha002;
m[13'd3918]=16'h4be1;
m[13'd3919]=16'h0408;
m[13'd3920]=16'h0009;
m[13'd3921]=16'h4907;
m[13'd3922]=16'h001b;
m[13'd3923]=16'h8009;
m[13'd3924]=16'h0010;
m[13'd3925]=16'h000a;
m[13'd3926]=16'h0015;
m[13'd3927]=16'h090c;
m[13'd3928]=16'h0009;
m[13'd3929]=16'h080d;
m[13'd3930]=16'h0007;
m[13'd3931]=16'h000b;
m[13'd3932]=16'h0009;
m[13'd3933]=16'h110b;
m[13'd3934]=16'h00c6;
m[13'd3935]=16'h0601;
m[13'd3936]=16'h0009;
m[13'd3937]=16'h6c00;
m[13'd3938]=16'h0018;
m[13'd3939]=16'h4104;
m[13'd3940]=16'h0025;
m[13'd3941]=16'h4004;
m[13'd3942]=16'h004e;
m[13'd3943]=16'h0003;
m[13'd3944]=16'h0009;
m[13'd3945]=16'hb002;
m[13'd3946]=16'h4a92;
m[13'd3947]=16'h810b;
m[13'd3948]=16'h003b;
m[13'd3949]=16'h0a08;
m[13'd3950]=16'h0009;
m[13'd3951]=16'hcd07;
m[13'd3952]=16'h0089;
m[13'd3953]=16'h0601;
m[13'd3954]=16'h0009;
m[13'd3955]=16'h6c00;
m[13'd3956]=16'h0018;
m[13'd3957]=16'h4104;
m[13'd3958]=16'h0025;
m[13'd3959]=16'h4004;
m[13'd3960]=16'h004e;
m[13'd3961]=16'h0003;
m[13'd3962]=16'h0009;
m[13'd3963]=16'hc002;
m[13'd3964]=16'h4b5d;
m[13'd3965]=16'h110b;
m[13'd3966]=16'h003b;
m[13'd3967]=16'h1108;
m[13'd3968]=16'h0009;
m[13'd3969]=16'h2507;
m[13'd3970]=16'h0089;
m[13'd3971]=16'h0601;
m[13'd3972]=16'h0009;
m[13'd3973]=16'h6c00;
m[13'd3974]=16'h0018;
m[13'd3975]=16'h4104;
m[13'd3976]=16'h0025;
m[13'd3977]=16'h4004;
m[13'd3978]=16'h004e;
m[13'd3979]=16'h0003;
m[13'd3980]=16'h0009;
m[13'd3981]=16'hd002;
m[13'd3982]=16'h4b60;
m[13'd3983]=16'h110b;
m[13'd3984]=16'h003b;
m[13'd3985]=16'h0d08;
m[13'd3986]=16'h0009;
m[13'd3987]=16'h9c07;
m[13'd3988]=16'h0089;
m[13'd3989]=16'h0601;
m[13'd3990]=16'h0009;
m[13'd3991]=16'h6c00;
m[13'd3992]=16'h0018;
m[13'd3993]=16'h4104;
m[13'd3994]=16'h0025;
m[13'd3995]=16'h4004;
m[13'd3996]=16'h004e;
m[13'd3997]=16'h0003;
m[13'd3998]=16'h0009;
m[13'd3999]=16'he002;
m[13'd4000]=16'h4b5d;
m[13'd4001]=16'h100b;
m[13'd4002]=16'h003b;
m[13'd4003]=16'h0a08;
m[13'd4004]=16'h0009;
m[13'd4005]=16'hcd07;
m[13'd4006]=16'h0089;
m[13'd4007]=16'h0601;
m[13'd4008]=16'h0009;
m[13'd4009]=16'h6c00;
m[13'd4010]=16'h0018;
m[13'd4011]=16'h4104;
m[13'd4012]=16'h0025;
m[13'd4013]=16'h4004;
m[13'd4014]=16'h004e;
m[13'd4015]=16'h0003;
m[13'd4016]=16'h0009;
m[13'd4017]=16'hf002;
m[13'd4018]=16'h4b5d;
m[13'd4019]=16'h100b;
m[13'd4020]=16'h003b;
m[13'd4021]=16'h0908;
m[13'd4022]=16'h0009;
m[13'd4023]=16'h9f07;
m[13'd4024]=16'h0089;
m[13'd4025]=16'h0601;
m[13'd4026]=16'h0009;
m[13'd4027]=16'h6c00;
m[13'd4028]=16'h0018;
m[13'd4029]=16'h4104;
m[13'd4030]=16'h0025;
m[13'd4031]=16'h4004;
m[13'd4032]=16'h004e;
m[13'd4033]=16'h0103;
m[13'd4034]=16'h0009;
m[13'd4035]=16'h0002;
m[13'd4036]=16'h4bd2;
m[13'd4037]=16'h0308;
m[13'd4038]=16'h0009;
m[13'd4039]=16'hd207;
m[13'd4040]=16'h001b;
m[13'd4041]=16'h8009;
m[13'd4042]=16'h0010;
m[13'd4043]=16'h000a;
m[13'd4044]=16'h0015;
m[13'd4045]=16'h090c;
m[13'd4046]=16'h0009;
m[13'd4047]=16'h080d;
m[13'd4048]=16'h0007;
m[13'd4049]=16'h000b;
m[13'd4050]=16'h0009;
m[13'd4051]=16'h110b;
m[13'd4052]=16'h015a;
m[13'd4053]=16'h0501;
m[13'd4054]=16'h0009;
m[13'd4055]=16'hb900;
m[13'd4056]=16'h001b;
m[13'd4057]=16'h4002;
m[13'd4058]=16'h0010;
m[13'd4059]=16'h0003;
m[13'd4060]=16'h0016;
m[13'd4061]=16'h0905;
m[13'd4062]=16'h000a;
m[13'd4063]=16'h0906;
m[13'd4064]=16'h0007;
m[13'd4065]=16'h0004;
m[13'd4066]=16'h000a;
m[13'd4067]=16'h4104;
m[13'd4068]=16'h008d;
m[13'd4069]=16'h0003;
m[13'd4070]=16'h0009;
m[13'd4071]=16'h5002;
m[13'd4072]=16'h499f;
m[13'd4073]=16'h810b;
m[13'd4074]=16'h003b;
m[13'd4075]=16'h0908;
m[13'd4076]=16'h0009;
m[13'd4077]=16'h9f07;
m[13'd4078]=16'h006a;
m[13'd4079]=16'h4801;
m[13'd4080]=16'h0007;
m[13'd4081]=16'h0000;
m[13'd4082]=16'h000e;
m[13'd4083]=16'h8104;
m[13'd4084]=16'h0058;
m[13'd4085]=16'h0003;
m[13'd4086]=16'h0009;
m[13'd4087]=16'h6002;
m[13'd4088]=16'h4ba2;
m[13'd4089]=16'h110b;
m[13'd4090]=16'h003b;
m[13'd4091]=16'h0f08;
m[13'd4092]=16'h0009;
m[13'd4093]=16'h4607;
m[13'd4094]=16'h0089;
m[13'd4095]=16'h0501;
m[13'd4096]=16'h0009;
m[13'd4097]=16'hb900;
m[13'd4098]=16'h0018;
m[13'd4099]=16'h4104;
m[13'd4100]=16'h0058;
m[13'd4101]=16'h0003;
m[13'd4102]=16'h0009;
m[13'd4103]=16'h7002;
m[13'd4104]=16'h4b7b;
m[13'd4105]=16'h110b;
m[13'd4106]=16'h003b;
m[13'd4107]=16'h0c08;
m[13'd4108]=16'h0009;
m[13'd4109]=16'h2007;
m[13'd4110]=16'h0089;
m[13'd4111]=16'h0501;
m[13'd4112]=16'h0009;
m[13'd4113]=16'hb900;
m[13'd4114]=16'h0018;
m[13'd4115]=16'h4104;
m[13'd4116]=16'h0058;
m[13'd4117]=16'h0003;
m[13'd4118]=16'h0009;
m[13'd4119]=16'h8002;
m[13'd4120]=16'h4b78;
m[13'd4121]=16'h100b;
m[13'd4122]=16'h003b;
m[13'd4123]=16'h0908;
m[13'd4124]=16'h0009;
m[13'd4125]=16'h9f07;
m[13'd4126]=16'h0089;
m[13'd4127]=16'h0501;
m[13'd4128]=16'h0009;
m[13'd4129]=16'hb900;
m[13'd4130]=16'h0018;
m[13'd4131]=16'h4104;
m[13'd4132]=16'h0058;
m[13'd4133]=16'h0003;
m[13'd4134]=16'h0009;
m[13'd4135]=16'h9002;
m[13'd4136]=16'h4b78;
m[13'd4137]=16'h100b;
m[13'd4138]=16'h003b;
m[13'd4139]=16'h0808;
m[13'd4140]=16'h0009;
m[13'd4141]=16'h9307;
m[13'd4142]=16'h0089;
m[13'd4143]=16'h0501;
m[13'd4144]=16'h0009;
m[13'd4145]=16'hb900;
m[13'd4146]=16'h0018;
m[13'd4147]=16'h4104;
m[13'd4148]=16'h0058;
m[13'd4149]=16'h0003;
m[13'd4150]=16'h0009;
m[13'd4151]=16'ha002;
m[13'd4152]=16'h4bfa;
m[13'd4153]=16'h0308;
m[13'd4154]=16'h0009;
m[13'd4155]=16'h6707;
m[13'd4156]=16'h001b;
m[13'd4157]=16'h8009;
m[13'd4158]=16'h0010;
m[13'd4159]=16'h000a;
m[13'd4160]=16'h0015;
m[13'd4161]=16'h090c;
m[13'd4162]=16'h0009;
m[13'd4163]=16'h080d;
m[13'd4164]=16'h0007;
m[13'd4165]=16'h000b;
m[13'd4166]=16'h0009;
m[13'd4167]=16'h110b;
m[13'd4168]=16'h0155;
m[13'd4169]=16'h0601;
m[13'd4170]=16'h0009;
m[13'd4171]=16'h6c00;
m[13'd4172]=16'h001b;
m[13'd4173]=16'h4002;
m[13'd4174]=16'h0010;
m[13'd4175]=16'h0003;
m[13'd4176]=16'h0016;
m[13'd4177]=16'h0905;
m[13'd4178]=16'h000a;
m[13'd4179]=16'h0906;
m[13'd4180]=16'h0007;
m[13'd4181]=16'h0004;
m[13'd4182]=16'h000a;
m[13'd4183]=16'h4104;
m[13'd4184]=16'h008d;
m[13'd4185]=16'h0003;
m[13'd4186]=16'h0009;
m[13'd4187]=16'h5002;
m[13'd4188]=16'h4996;
m[13'd4189]=16'h810b;
m[13'd4190]=16'h003b;
m[13'd4191]=16'h0808;
m[13'd4192]=16'h0009;
m[13'd4193]=16'h9307;
m[13'd4194]=16'h0072;
m[13'd4195]=16'h4801;
m[13'd4196]=16'h0007;
m[13'd4197]=16'h0000;
m[13'd4198]=16'h000e;
m[13'd4199]=16'h8104;
m[13'd4200]=16'h0058;
m[13'd4201]=16'h0003;
m[13'd4202]=16'h0009;
m[13'd4203]=16'h6002;
m[13'd4204]=16'h4b9c;
m[13'd4205]=16'h110b;
m[13'd4206]=16'h003b;
m[13'd4207]=16'h0d08;
m[13'd4208]=16'h0009;
m[13'd4209]=16'h9c07;
m[13'd4210]=16'h0091;
m[13'd4211]=16'h0601;
m[13'd4212]=16'h0009;
m[13'd4213]=16'h6c00;
m[13'd4214]=16'h0018;
m[13'd4215]=16'h4104;
m[13'd4216]=16'h0058;
m[13'd4217]=16'h0003;
m[13'd4218]=16'h0009;
m[13'd4219]=16'h7002;
m[13'd4220]=16'h4b72;
m[13'd4221]=16'h110b;
m[13'd4222]=16'h003b;
m[13'd4223]=16'h0a08;
m[13'd4224]=16'h0009;
m[13'd4225]=16'hcd07;
m[13'd4226]=16'h0091;
m[13'd4227]=16'h0601;
m[13'd4228]=16'h0009;
m[13'd4229]=16'h6c00;
m[13'd4230]=16'h0018;
m[13'd4231]=16'h4104;
m[13'd4232]=16'h0058;
m[13'd4233]=16'h0003;
m[13'd4234]=16'h0009;
m[13'd4235]=16'h8002;
m[13'd4236]=16'h4b6f;
m[13'd4237]=16'h100b;
m[13'd4238]=16'h003b;
m[13'd4239]=16'h0808;
m[13'd4240]=16'h0009;
m[13'd4241]=16'h9307;
m[13'd4242]=16'h0091;
m[13'd4243]=16'h0601;
m[13'd4244]=16'h0009;
m[13'd4245]=16'h6c00;
m[13'd4246]=16'h0018;
m[13'd4247]=16'h4104;
m[13'd4248]=16'h0058;
m[13'd4249]=16'h0003;
m[13'd4250]=16'h0009;
m[13'd4251]=16'h9002;
m[13'd4252]=16'h4b72;
m[13'd4253]=16'h100b;
m[13'd4254]=16'h003b;
m[13'd4255]=16'h0708;
m[13'd4256]=16'h0009;
m[13'd4257]=16'ha307;
m[13'd4258]=16'h0091;
m[13'd4259]=16'h0601;
m[13'd4260]=16'h0009;
m[13'd4261]=16'h6c00;
m[13'd4262]=16'h0018;
m[13'd4263]=16'h4104;
m[13'd4264]=16'h0058;
m[13'd4265]=16'h0003;
m[13'd4266]=16'h0009;
m[13'd4267]=16'ha002;
m[13'd4268]=16'h4b82;
m[13'd4269]=16'h100b;
m[13'd4270]=16'h003b;
m[13'd4271]=16'h0608;
m[13'd4272]=16'h0009;
m[13'd4273]=16'hce07;
m[13'd4274]=16'h0024;
m[13'd4275]=16'h100b;
m[13'd4276]=16'h010e;
m[13'd4277]=16'h0601;
m[13'd4278]=16'h0009;
m[13'd4279]=16'hce00;
m[13'd4280]=16'h001b;
m[13'd4281]=16'h4002;
m[13'd4282]=16'h0010;
m[13'd4283]=16'h0003;
m[13'd4284]=16'h0016;
m[13'd4285]=16'h0905;
m[13'd4286]=16'h000a;
m[13'd4287]=16'h0906;
m[13'd4288]=16'h0007;
m[13'd4289]=16'h0004;
m[13'd4290]=16'h000a;
m[13'd4291]=16'h4104;
m[13'd4292]=16'h008d;
m[13'd4293]=16'h0003;
m[13'd4294]=16'h0009;
m[13'd4295]=16'h5002;
m[13'd4296]=16'h4a47;
m[13'd4297]=16'h100b;
m[13'd4298]=16'h003b;
m[13'd4299]=16'h0608;
m[13'd4300]=16'h0009;
m[13'd4301]=16'h1007;
m[13'd4302]=16'h0024;
m[13'd4303]=16'h100b;
m[13'd4304]=16'h0060;
m[13'd4305]=16'h4801;
m[13'd4306]=16'h0007;
m[13'd4307]=16'h0000;
m[13'd4308]=16'h000e;
m[13'd4309]=16'h8104;
m[13'd4310]=16'h0058;
m[13'd4311]=16'h0003;
m[13'd4312]=16'h0009;
m[13'd4313]=16'h6002;
m[13'd4314]=16'h4b8a;
m[13'd4315]=16'h100b;
m[13'd4316]=16'h003a;
m[13'd4317]=16'h0508;
m[13'd4318]=16'h0009;
m[13'd4319]=16'h6707;
m[13'd4320]=16'h0024;
m[13'd4321]=16'h100b;
m[13'd4322]=16'h007f;
m[13'd4323]=16'h0601;
m[13'd4324]=16'h0009;
m[13'd4325]=16'hce00;
m[13'd4326]=16'h0018;
m[13'd4327]=16'h4104;
m[13'd4328]=16'h0058;
m[13'd4329]=16'h0003;
m[13'd4330]=16'h0009;
m[13'd4331]=16'h7002;
m[13'd4332]=16'h4b60;
m[13'd4333]=16'h100b;
m[13'd4334]=16'h003a;
m[13'd4335]=16'h0408;
m[13'd4336]=16'h0009;
m[13'd4337]=16'hd007;
m[13'd4338]=16'h0024;
m[13'd4339]=16'h100b;
m[13'd4340]=16'h007f;
m[13'd4341]=16'h0601;
m[13'd4342]=16'h0009;
m[13'd4343]=16'hce00;
m[13'd4344]=16'h0018;
m[13'd4345]=16'h4104;
m[13'd4346]=16'h0058;
m[13'd4347]=16'h0003;
m[13'd4348]=16'h0009;
m[13'd4349]=16'h8002;
m[13'd4350]=16'h4b60;
m[13'd4351]=16'h100b;
m[13'd4352]=16'h003a;
m[13'd4353]=16'h0408;
m[13'd4354]=16'h0009;
m[13'd4355]=16'h4907;
m[13'd4356]=16'h0024;
m[13'd4357]=16'h100b;
m[13'd4358]=16'h007f;
m[13'd4359]=16'h0601;
m[13'd4360]=16'h0009;
m[13'd4361]=16'hce00;
m[13'd4362]=16'h0018;
m[13'd4363]=16'h4104;
m[13'd4364]=16'h0058;
m[13'd4365]=16'h0003;
m[13'd4366]=16'h0009;
m[13'd4367]=16'h9002;
m[13'd4368]=16'h4b60;
m[13'd4369]=16'h100b;
m[13'd4370]=16'h003a;
m[13'd4371]=16'h0308;
m[13'd4372]=16'h0009;
m[13'd4373]=16'hd207;
m[13'd4374]=16'h0024;
m[13'd4375]=16'h100b;
m[13'd4376]=16'h007f;
m[13'd4377]=16'h0601;
m[13'd4378]=16'h0009;
m[13'd4379]=16'hce00;
m[13'd4380]=16'h0018;
m[13'd4381]=16'h4104;
m[13'd4382]=16'h0058;
m[13'd4383]=16'h0003;
m[13'd4384]=16'h0009;
m[13'd4385]=16'ha002;
m[13'd4386]=16'h4bff;
m[13'd4387]=16'h000f;
m[13'd4388]=16'h0009;
m[13'd4389]=16'h000e;
m[13'd4390]=16'h001b;
m[13'd4391]=16'h0010;
m[13'd4392]=16'h0010;
m[13'd4393]=16'h0011;
m[13'd4394]=16'h0015;
m[13'd4395]=16'h0013;
m[13'd4396]=16'h0009;
m[13'd4397]=16'h0014;
m[13'd4398]=16'h0007;
m[13'd4399]=16'h0012;
m[13'd4400]=16'h0009;
m[13'd4401]=16'h4012;
m[13'd4402]=16'h01e0;
m[13'd4403]=16'h0708;
m[13'd4404]=16'h0009;
m[13'd4405]=16'h3507;
m[13'd4406]=16'h001b;
m[13'd4407]=16'h4009;
m[13'd4408]=16'h0010;
m[13'd4409]=16'h000a;
m[13'd4410]=16'h0016;
m[13'd4411]=16'h090c;
m[13'd4412]=16'h000a;
m[13'd4413]=16'h090d;
m[13'd4414]=16'h0007;
m[13'd4415]=16'h000b;
m[13'd4416]=16'h000a;
m[13'd4417]=16'h410b;
m[13'd4418]=16'h0095;
m[13'd4419]=16'h000a;
m[13'd4420]=16'h0009;
m[13'd4421]=16'h5009;
m[13'd4422]=16'h0176;
m[13'd4423]=16'h0301;
m[13'd4424]=16'h0009;
m[13'd4425]=16'h9b00;
m[13'd4426]=16'h001b;
m[13'd4427]=16'h4002;
m[13'd4428]=16'h0010;
m[13'd4429]=16'h0003;
m[13'd4430]=16'h0016;
m[13'd4431]=16'h0905;
m[13'd4432]=16'h000a;
m[13'd4433]=16'h0906;
m[13'd4434]=16'h0007;
m[13'd4435]=16'h0004;
m[13'd4436]=16'h000a;
m[13'd4437]=16'h4104;
m[13'd4438]=16'h0095;
m[13'd4439]=16'h0003;
m[13'd4440]=16'h0009;
m[13'd4441]=16'h5002;
m[13'd4442]=16'h46a5;
m[13'd4443]=16'h000a;
m[13'd4444]=16'h0009;
m[13'd4445]=16'h6009;
m[13'd4446]=16'h0055;
m[13'd4447]=16'h4801;
m[13'd4448]=16'h0007;
m[13'd4449]=16'h0000;
m[13'd4450]=16'h000e;
m[13'd4451]=16'h8104;
m[13'd4452]=16'h0060;
m[13'd4453]=16'h0003;
m[13'd4454]=16'h0009;
m[13'd4455]=16'h6002;
m[13'd4456]=16'h4bed;
m[13'd4457]=16'h000a;
m[13'd4458]=16'h0009;
m[13'd4459]=16'h7009;
m[13'd4460]=16'h0073;
m[13'd4461]=16'h0301;
m[13'd4462]=16'h0009;
m[13'd4463]=16'h9b00;
m[13'd4464]=16'h0018;
m[13'd4465]=16'h4104;
m[13'd4466]=16'h0060;
m[13'd4467]=16'h0003;
m[13'd4468]=16'h0009;
m[13'd4469]=16'h7002;
m[13'd4470]=16'h4bc3;
m[13'd4471]=16'h000a;
m[13'd4472]=16'h0009;
m[13'd4473]=16'h8009;
m[13'd4474]=16'h0073;
m[13'd4475]=16'h0301;
m[13'd4476]=16'h0009;
m[13'd4477]=16'h9b00;
m[13'd4478]=16'h0018;
m[13'd4479]=16'h4104;
m[13'd4480]=16'h0060;
m[13'd4481]=16'h0003;
m[13'd4482]=16'h0009;
m[13'd4483]=16'h8002;
m[13'd4484]=16'h4bc0;
m[13'd4485]=16'h000a;
m[13'd4486]=16'h0009;
m[13'd4487]=16'h9009;
m[13'd4488]=16'h0073;
m[13'd4489]=16'h0301;
m[13'd4490]=16'h0009;
m[13'd4491]=16'h9b00;
m[13'd4492]=16'h0018;
m[13'd4493]=16'h4104;
m[13'd4494]=16'h0060;
m[13'd4495]=16'h0003;
m[13'd4496]=16'h0009;
m[13'd4497]=16'h9002;
m[13'd4498]=16'h4bc3;
m[13'd4499]=16'h000a;
m[13'd4500]=16'h0009;
m[13'd4501]=16'ha009;
m[13'd4502]=16'h0073;
m[13'd4503]=16'h0301;
m[13'd4504]=16'h0009;
m[13'd4505]=16'h9b00;
m[13'd4506]=16'h0018;
m[13'd4507]=16'h4104;
m[13'd4508]=16'h0060;
m[13'd4509]=16'h0003;
m[13'd4510]=16'h0009;
m[13'd4511]=16'ha002;
m[13'd4512]=16'h4bd3;
m[13'd4513]=16'h000a;
m[13'd4514]=16'h0009;
m[13'd4515]=16'hb009;
m[13'd4516]=16'h007b;
m[13'd4517]=16'h0301;
m[13'd4518]=16'h0009;
m[13'd4519]=16'h9b00;
m[13'd4520]=16'h0018;
m[13'd4521]=16'h4104;
m[13'd4522]=16'h0025;
m[13'd4523]=16'h4004;
m[13'd4524]=16'h004e;
m[13'd4525]=16'h0003;
m[13'd4526]=16'h0009;
m[13'd4527]=16'hb002;
m[13'd4528]=16'h4b97;
m[13'd4529]=16'h000a;
m[13'd4530]=16'h0009;
m[13'd4531]=16'hc009;
m[13'd4532]=16'h0073;
m[13'd4533]=16'h0301;
m[13'd4534]=16'h0009;
m[13'd4535]=16'h9b00;
m[13'd4536]=16'h0018;
m[13'd4537]=16'h4104;
m[13'd4538]=16'h0025;
m[13'd4539]=16'h4004;
m[13'd4540]=16'h004e;
m[13'd4541]=16'h0003;
m[13'd4542]=16'h0009;
m[13'd4543]=16'hc002;
m[13'd4544]=16'h4bae;
m[13'd4545]=16'h000a;
m[13'd4546]=16'h0009;
m[13'd4547]=16'hd009;
m[13'd4548]=16'h0073;
m[13'd4549]=16'h0301;
m[13'd4550]=16'h0009;
m[13'd4551]=16'h9b00;
m[13'd4552]=16'h0018;
m[13'd4553]=16'h4104;
m[13'd4554]=16'h0025;
m[13'd4555]=16'h4004;
m[13'd4556]=16'h004e;
m[13'd4557]=16'h0003;
m[13'd4558]=16'h0009;
m[13'd4559]=16'hd002;
m[13'd4560]=16'h4bae;
m[13'd4561]=16'h000a;
m[13'd4562]=16'h0009;
m[13'd4563]=16'he009;
m[13'd4564]=16'h0073;
m[13'd4565]=16'h0301;
m[13'd4566]=16'h0009;
m[13'd4567]=16'h9b00;
m[13'd4568]=16'h0018;
m[13'd4569]=16'h4104;
m[13'd4570]=16'h0025;
m[13'd4571]=16'h4004;
m[13'd4572]=16'h004e;
m[13'd4573]=16'h0003;
m[13'd4574]=16'h0009;
m[13'd4575]=16'he002;
m[13'd4576]=16'h4bb1;
m[13'd4577]=16'h000a;
m[13'd4578]=16'h0009;
m[13'd4579]=16'hf009;
m[13'd4580]=16'h0073;
m[13'd4581]=16'h0301;
m[13'd4582]=16'h0009;
m[13'd4583]=16'h9b00;
m[13'd4584]=16'h0018;
m[13'd4585]=16'h4104;
m[13'd4586]=16'h0025;
m[13'd4587]=16'h4004;
m[13'd4588]=16'h004e;
m[13'd4589]=16'h0003;
m[13'd4590]=16'h0009;
m[13'd4591]=16'hf002;
m[13'd4592]=16'h4bae;
m[13'd4593]=16'h010a;
m[13'd4594]=16'h0009;
m[13'd4595]=16'h0009;
m[13'd4596]=16'h0073;
m[13'd4597]=16'h0301;
m[13'd4598]=16'h0009;
m[13'd4599]=16'h9b00;
m[13'd4600]=16'h0018;
m[13'd4601]=16'h4104;
m[13'd4602]=16'h0025;
m[13'd4603]=16'h4004;
m[13'd4604]=16'h004e;
m[13'd4605]=16'h0103;
m[13'd4606]=16'h0009;
m[13'd4607]=16'h0002;
m[13'd4608]=16'h4b83;
m[13'd4609]=16'h400b;
m[13'd4610]=16'h004e;
m[13'd4611]=16'h010a;
m[13'd4612]=16'h0009;
m[13'd4613]=16'h1009;
m[13'd4614]=16'h0102;
m[13'd4615]=16'h0301;
m[13'd4616]=16'h0009;
m[13'd4617]=16'h9b00;
m[13'd4618]=16'h001b;
m[13'd4619]=16'h4002;
m[13'd4620]=16'h0010;
m[13'd4621]=16'h0003;
m[13'd4622]=16'h0016;
m[13'd4623]=16'h0905;
m[13'd4624]=16'h000a;
m[13'd4625]=16'h0906;
m[13'd4626]=16'h0007;
m[13'd4627]=16'h0004;
m[13'd4628]=16'h000a;
m[13'd4629]=16'h4104;
m[13'd4630]=16'h0095;
m[13'd4631]=16'h0003;
m[13'd4632]=16'h0009;
m[13'd4633]=16'h5002;
m[13'd4634]=16'h4a5d;
m[13'd4635]=16'h400b;
m[13'd4636]=16'h004e;
m[13'd4637]=16'h010a;
m[13'd4638]=16'h0009;
m[13'd4639]=16'h2009;
m[13'd4640]=16'h0055;
m[13'd4641]=16'h4801;
m[13'd4642]=16'h0007;
m[13'd4643]=16'h0000;
m[13'd4644]=16'h000e;
m[13'd4645]=16'h8104;
m[13'd4646]=16'h0060;
m[13'd4647]=16'h0003;
m[13'd4648]=16'h0009;
m[13'd4649]=16'h6002;
m[13'd4650]=16'h4b9d;
m[13'd4651]=16'h400b;
m[13'd4652]=16'h004e;
m[13'd4653]=16'h010a;
m[13'd4654]=16'h0009;
m[13'd4655]=16'h3009;
m[13'd4656]=16'h0073;
m[13'd4657]=16'h0301;
m[13'd4658]=16'h0009;
m[13'd4659]=16'h9b00;
m[13'd4660]=16'h0018;
m[13'd4661]=16'h4104;
m[13'd4662]=16'h0060;
m[13'd4663]=16'h0003;
m[13'd4664]=16'h0009;
m[13'd4665]=16'h7002;
m[13'd4666]=16'h4b76;
m[13'd4667]=16'h400b;
m[13'd4668]=16'h004e;
m[13'd4669]=16'h010a;
m[13'd4670]=16'h0009;
m[13'd4671]=16'h4009;
m[13'd4672]=16'h0073;
m[13'd4673]=16'h0301;
m[13'd4674]=16'h0009;
m[13'd4675]=16'h9b00;
m[13'd4676]=16'h0018;
m[13'd4677]=16'h4104;
m[13'd4678]=16'h0060;
m[13'd4679]=16'h0003;
m[13'd4680]=16'h0009;
m[13'd4681]=16'h8002;
m[13'd4682]=16'h4b73;
m[13'd4683]=16'h400b;
m[13'd4684]=16'h004e;
m[13'd4685]=16'h010a;
m[13'd4686]=16'h0009;
m[13'd4687]=16'h5009;
m[13'd4688]=16'h0073;
m[13'd4689]=16'h0301;
m[13'd4690]=16'h0009;
m[13'd4691]=16'h9b00;
m[13'd4692]=16'h0018;
m[13'd4693]=16'h4104;
m[13'd4694]=16'h0060;
m[13'd4695]=16'h0003;
m[13'd4696]=16'h0009;
m[13'd4697]=16'h9002;
m[13'd4698]=16'h4b73;
m[13'd4699]=16'h400b;
m[13'd4700]=16'h004e;
m[13'd4701]=16'h010a;
m[13'd4702]=16'h0009;
m[13'd4703]=16'h6009;
m[13'd4704]=16'h0073;
m[13'd4705]=16'h0301;
m[13'd4706]=16'h0009;
m[13'd4707]=16'h9b00;
m[13'd4708]=16'h0018;
m[13'd4709]=16'h4104;
m[13'd4710]=16'h0060;
m[13'd4711]=16'h0003;
m[13'd4712]=16'h0009;
m[13'd4713]=16'ha002;
m[13'd4714]=16'h4bc1;
m[13'd4715]=16'h010a;
m[13'd4716]=16'h0009;
m[13'd4717]=16'h7009;
m[13'd4718]=16'h007b;
m[13'd4719]=16'h0301;
m[13'd4720]=16'h0009;
m[13'd4721]=16'h9b00;
m[13'd4722]=16'h0018;
m[13'd4723]=16'h4104;
m[13'd4724]=16'h0025;
m[13'd4725]=16'h4004;
m[13'd4726]=16'h004e;
m[13'd4727]=16'h0003;
m[13'd4728]=16'h0009;
m[13'd4729]=16'hb002;
m[13'd4730]=16'h4b97;
m[13'd4731]=16'h010a;
m[13'd4732]=16'h0009;
m[13'd4733]=16'h8009;
m[13'd4734]=16'h0073;
m[13'd4735]=16'h0301;
m[13'd4736]=16'h0009;
m[13'd4737]=16'h9b00;
m[13'd4738]=16'h0018;
m[13'd4739]=16'h4104;
m[13'd4740]=16'h0025;
m[13'd4741]=16'h4004;
m[13'd4742]=16'h004e;
m[13'd4743]=16'h0003;
m[13'd4744]=16'h0009;
m[13'd4745]=16'hc002;
m[13'd4746]=16'h4bae;
m[13'd4747]=16'h010a;
m[13'd4748]=16'h0009;
m[13'd4749]=16'h9009;
m[13'd4750]=16'h0073;
m[13'd4751]=16'h0301;
m[13'd4752]=16'h0009;
m[13'd4753]=16'h9b00;
m[13'd4754]=16'h0018;
m[13'd4755]=16'h4104;
m[13'd4756]=16'h0025;
m[13'd4757]=16'h4004;
m[13'd4758]=16'h004e;
m[13'd4759]=16'h0003;
m[13'd4760]=16'h0009;
m[13'd4761]=16'hd002;
m[13'd4762]=16'h4bae;
m[13'd4763]=16'h010a;
m[13'd4764]=16'h0009;
m[13'd4765]=16'ha009;
m[13'd4766]=16'h0073;
m[13'd4767]=16'h0301;
m[13'd4768]=16'h0009;
m[13'd4769]=16'h9b00;
m[13'd4770]=16'h0018;
m[13'd4771]=16'h4104;
m[13'd4772]=16'h0025;
m[13'd4773]=16'h4004;
m[13'd4774]=16'h004e;
m[13'd4775]=16'h0003;
m[13'd4776]=16'h0009;
m[13'd4777]=16'he002;
m[13'd4778]=16'h4bb1;
m[13'd4779]=16'h010a;
m[13'd4780]=16'h0009;
m[13'd4781]=16'hb009;
m[13'd4782]=16'h0073;
m[13'd4783]=16'h0301;
m[13'd4784]=16'h0009;
m[13'd4785]=16'h9b00;
m[13'd4786]=16'h0018;
m[13'd4787]=16'h4104;
m[13'd4788]=16'h0025;
m[13'd4789]=16'h4004;
m[13'd4790]=16'h004e;
m[13'd4791]=16'h0003;
m[13'd4792]=16'h0009;
m[13'd4793]=16'hf002;
m[13'd4794]=16'h4bae;
m[13'd4795]=16'h010a;
m[13'd4796]=16'h0009;
m[13'd4797]=16'hc009;
m[13'd4798]=16'h0073;
m[13'd4799]=16'h0301;
m[13'd4800]=16'h0009;
m[13'd4801]=16'h9b00;
m[13'd4802]=16'h0018;
m[13'd4803]=16'h4104;
m[13'd4804]=16'h0025;
m[13'd4805]=16'h4004;
m[13'd4806]=16'h004e;
m[13'd4807]=16'h0103;
m[13'd4808]=16'h0009;
m[13'd4809]=16'h0002;
m[13'd4810]=16'h4c0b;
m[13'd4811]=16'h0108;
m[13'd4812]=16'h0009;
m[13'd4813]=16'h2307;
m[13'd4814]=16'h001b;
m[13'd4815]=16'h4009;
m[13'd4816]=16'h0010;
m[13'd4817]=16'h000a;
m[13'd4818]=16'h0016;
m[13'd4819]=16'h090c;
m[13'd4820]=16'h000a;
m[13'd4821]=16'h090d;
m[13'd4822]=16'h0007;
m[13'd4823]=16'h000b;
m[13'd4824]=16'h000a;
m[13'd4825]=16'h410b;
m[13'd4826]=16'h0095;
m[13'd4827]=16'h000a;
m[13'd4828]=16'h0009;
m[13'd4829]=16'h5009;
m[13'd4830]=16'h010f;
m[13'd4831]=16'h0301;
m[13'd4832]=16'h0009;
m[13'd4833]=16'h9b00;
m[13'd4834]=16'h001b;
m[13'd4835]=16'h4002;
m[13'd4836]=16'h0010;
m[13'd4837]=16'h0003;
m[13'd4838]=16'h0016;
m[13'd4839]=16'h0905;
m[13'd4840]=16'h000a;
m[13'd4841]=16'h0906;
m[13'd4842]=16'h0007;
m[13'd4843]=16'h0004;
m[13'd4844]=16'h000a;
m[13'd4845]=16'h4104;
m[13'd4846]=16'h008d;
m[13'd4847]=16'h0003;
m[13'd4848]=16'h0009;
m[13'd4849]=16'h5002;
m[13'd4850]=16'h4927;
m[13'd4851]=16'h810b;
m[13'd4852]=16'h002b;
m[13'd4853]=16'h3108;
m[13'd4854]=16'h0007;
m[13'd4855]=16'h0007;
m[13'd4856]=16'h0060;
m[13'd4857]=16'h000a;
m[13'd4858]=16'h0009;
m[13'd4859]=16'h6009;
m[13'd4860]=16'h0055;
m[13'd4861]=16'h4801;
m[13'd4862]=16'h0007;
m[13'd4863]=16'h0000;
m[13'd4864]=16'h000e;
m[13'd4865]=16'h8104;
m[13'd4866]=16'h0058;
m[13'd4867]=16'h0003;
m[13'd4868]=16'h0009;
m[13'd4869]=16'h6002;
m[13'd4870]=16'h4b60;
m[13'd4871]=16'h110b;
m[13'd4872]=16'h002b;
m[13'd4873]=16'h1108;
m[13'd4874]=16'h0007;
m[13'd4875]=16'h0007;
m[13'd4876]=16'h0060;
m[13'd4877]=16'h000a;
m[13'd4878]=16'h0009;
m[13'd4879]=16'h7009;
m[13'd4880]=16'h0073;
m[13'd4881]=16'h0301;
m[13'd4882]=16'h0009;
m[13'd4883]=16'h9b00;
m[13'd4884]=16'h0018;
m[13'd4885]=16'h4104;
m[13'd4886]=16'h0058;
m[13'd4887]=16'h0003;
m[13'd4888]=16'h0009;
m[13'd4889]=16'h7002;
m[13'd4890]=16'h4b39;
m[13'd4891]=16'h800b;
m[13'd4892]=16'h002b;
m[13'd4893]=16'h0808;
m[13'd4894]=16'h0007;
m[13'd4895]=16'h0007;
m[13'd4896]=16'h0060;
m[13'd4897]=16'h000a;
m[13'd4898]=16'h0009;
m[13'd4899]=16'h8009;
m[13'd4900]=16'h0073;
m[13'd4901]=16'h0301;
m[13'd4902]=16'h0009;
m[13'd4903]=16'h9b00;
m[13'd4904]=16'h0018;
m[13'd4905]=16'h4104;
m[13'd4906]=16'h0058;
m[13'd4907]=16'h0003;
m[13'd4908]=16'h0009;
m[13'd4909]=16'h8002;
m[13'd4910]=16'h4b39;
m[13'd4911]=16'h400b;
m[13'd4912]=16'h002b;
m[13'd4913]=16'h1608;
m[13'd4914]=16'h0007;
m[13'd4915]=16'h0007;
m[13'd4916]=16'h0060;
m[13'd4917]=16'h000a;
m[13'd4918]=16'h0009;
m[13'd4919]=16'h9009;
m[13'd4920]=16'h0073;
m[13'd4921]=16'h0301;
m[13'd4922]=16'h0009;
m[13'd4923]=16'h9b00;
m[13'd4924]=16'h0018;
m[13'd4925]=16'h4104;
m[13'd4926]=16'h0058;
m[13'd4927]=16'h0003;
m[13'd4928]=16'h0009;
m[13'd4929]=16'h9002;
m[13'd4930]=16'h4b36;
m[13'd4931]=16'h800b;
m[13'd4932]=16'h002b;
m[13'd4933]=16'h0508;
m[13'd4934]=16'h0007;
m[13'd4935]=16'h0007;
m[13'd4936]=16'h0060;
m[13'd4937]=16'h000a;
m[13'd4938]=16'h0009;
m[13'd4939]=16'ha009;
m[13'd4940]=16'h0073;
m[13'd4941]=16'h0301;
m[13'd4942]=16'h0009;
m[13'd4943]=16'h9b00;
m[13'd4944]=16'h0018;
m[13'd4945]=16'h4104;
m[13'd4946]=16'h0058;
m[13'd4947]=16'h0003;
m[13'd4948]=16'h0009;
m[13'd4949]=16'ha002;
m[13'd4950]=16'h4b49;
m[13'd4951]=16'h800b;
m[13'd4952]=16'h002b;
m[13'd4953]=16'h0408;
m[13'd4954]=16'h0007;
m[13'd4955]=16'h0007;
m[13'd4956]=16'h0025;
m[13'd4957]=16'h400b;
m[13'd4958]=16'h004e;
m[13'd4959]=16'h000a;
m[13'd4960]=16'h0009;
m[13'd4961]=16'hb009;
m[13'd4962]=16'h0102;
m[13'd4963]=16'h0401;
m[13'd4964]=16'h0009;
m[13'd4965]=16'h4900;
m[13'd4966]=16'h001b;
m[13'd4967]=16'h4002;
m[13'd4968]=16'h0010;
m[13'd4969]=16'h0003;
m[13'd4970]=16'h0016;
m[13'd4971]=16'h0905;
m[13'd4972]=16'h000a;
m[13'd4973]=16'h0906;
m[13'd4974]=16'h0007;
m[13'd4975]=16'h0004;
m[13'd4976]=16'h000a;
m[13'd4977]=16'h4104;
m[13'd4978]=16'h008d;
m[13'd4979]=16'h0003;
m[13'd4980]=16'h0009;
m[13'd4981]=16'h5002;
m[13'd4982]=16'h4a0e;
m[13'd4983]=16'h800b;
m[13'd4984]=16'h002b;
m[13'd4985]=16'h0308;
m[13'd4986]=16'h0007;
m[13'd4987]=16'h0007;
m[13'd4988]=16'h0025;
m[13'd4989]=16'h400b;
m[13'd4990]=16'h004e;
m[13'd4991]=16'h000a;
m[13'd4992]=16'h0009;
m[13'd4993]=16'hc009;
m[13'd4994]=16'h0055;
m[13'd4995]=16'h4801;
m[13'd4996]=16'h0007;
m[13'd4997]=16'h0000;
m[13'd4998]=16'h000e;
m[13'd4999]=16'h8104;
m[13'd5000]=16'h0058;
m[13'd5001]=16'h0003;
m[13'd5002]=16'h0009;
m[13'd5003]=16'h6002;
m[13'd5004]=16'h4b4e;
m[13'd5005]=16'h800b;
m[13'd5006]=16'h002b;
m[13'd5007]=16'h0308;
m[13'd5008]=16'h0007;
m[13'd5009]=16'h0007;
m[13'd5010]=16'h0025;
m[13'd5011]=16'h400b;
m[13'd5012]=16'h004e;
m[13'd5013]=16'h000a;
m[13'd5014]=16'h0009;
m[13'd5015]=16'hd009;
m[13'd5016]=16'h0073;
m[13'd5017]=16'h0401;
m[13'd5018]=16'h0009;
m[13'd5019]=16'h4900;
m[13'd5020]=16'h0018;
m[13'd5021]=16'h4104;
m[13'd5022]=16'h0058;
m[13'd5023]=16'h0003;
m[13'd5024]=16'h0009;
m[13'd5025]=16'h7002;
m[13'd5026]=16'h4b24;
m[13'd5027]=16'h100b;
m[13'd5028]=16'h002b;
m[13'd5029]=16'h1208;
m[13'd5030]=16'h0007;
m[13'd5031]=16'h0007;
m[13'd5032]=16'h0025;
m[13'd5033]=16'h400b;
m[13'd5034]=16'h004e;
m[13'd5035]=16'h000a;
m[13'd5036]=16'h0009;
m[13'd5037]=16'he009;
m[13'd5038]=16'h0073;
m[13'd5039]=16'h0401;
m[13'd5040]=16'h0009;
m[13'd5041]=16'h4900;
m[13'd5042]=16'h0018;
m[13'd5043]=16'h4104;
m[13'd5044]=16'h0058;
m[13'd5045]=16'h0003;
m[13'd5046]=16'h0009;
m[13'd5047]=16'h8002;
m[13'd5048]=16'h4b27;
m[13'd5049]=16'h100b;
m[13'd5050]=16'h002b;
m[13'd5051]=16'h1208;
m[13'd5052]=16'h0007;
m[13'd5053]=16'h0007;
m[13'd5054]=16'h0025;
m[13'd5055]=16'h400b;
m[13'd5056]=16'h004e;
m[13'd5057]=16'h000a;
m[13'd5058]=16'h0009;
m[13'd5059]=16'hf009;
m[13'd5060]=16'h0073;
m[13'd5061]=16'h0401;
m[13'd5062]=16'h0009;
m[13'd5063]=16'h4900;
m[13'd5064]=16'h0018;
m[13'd5065]=16'h4104;
m[13'd5066]=16'h0058;
m[13'd5067]=16'h0003;
m[13'd5068]=16'h0009;
m[13'd5069]=16'h9002;
m[13'd5070]=16'h4b24;
m[13'd5071]=16'h100b;
m[13'd5072]=16'h002b;
m[13'd5073]=16'h1108;
m[13'd5074]=16'h0007;
m[13'd5075]=16'h0007;
m[13'd5076]=16'h0025;
m[13'd5077]=16'h400b;
m[13'd5078]=16'h004e;
m[13'd5079]=16'h010a;
m[13'd5080]=16'h0009;
m[13'd5081]=16'h0009;
m[13'd5082]=16'h0073;
m[13'd5083]=16'h0401;
m[13'd5084]=16'h0009;
m[13'd5085]=16'h4900;
m[13'd5086]=16'h0018;
m[13'd5087]=16'h4104;
m[13'd5088]=16'h0058;
m[13'd5089]=16'h0003;
m[13'd5090]=16'h0009;
m[13'd5091]=16'ha002;
m[13'd5092]=16'h4bae;
m[13'd5093]=16'h0808;
m[13'd5094]=16'h0009;
m[13'd5095]=16'h9307;
m[13'd5096]=16'h001b;
m[13'd5097]=16'h4009;
m[13'd5098]=16'h0010;
m[13'd5099]=16'h000a;
m[13'd5100]=16'h0016;
m[13'd5101]=16'h090c;
m[13'd5102]=16'h000a;
m[13'd5103]=16'h090d;
m[13'd5104]=16'h0007;
m[13'd5105]=16'h000b;
m[13'd5106]=16'h000a;
m[13'd5107]=16'h410b;
m[13'd5108]=16'h0095;
m[13'd5109]=16'h000a;
m[13'd5110]=16'h0009;
m[13'd5111]=16'h5009;
m[13'd5112]=16'h010f;
m[13'd5113]=16'h0301;
m[13'd5114]=16'h0009;
m[13'd5115]=16'h9b00;
m[13'd5116]=16'h001b;
m[13'd5117]=16'h4002;
m[13'd5118]=16'h0010;
m[13'd5119]=16'h0003;
m[13'd5120]=16'h0016;
m[13'd5121]=16'h0905;
m[13'd5122]=16'h000a;
m[13'd5123]=16'h0906;
m[13'd5124]=16'h0007;
m[13'd5125]=16'h0004;
m[13'd5126]=16'h000a;
m[13'd5127]=16'h4104;
m[13'd5128]=16'h0095;
m[13'd5129]=16'h0003;
m[13'd5130]=16'h0009;
m[13'd5131]=16'h5002;
m[13'd5132]=16'h4963;
m[13'd5133]=16'h000a;
m[13'd5134]=16'h0009;
m[13'd5135]=16'h6009;
m[13'd5136]=16'h0055;
m[13'd5137]=16'h4801;
m[13'd5138]=16'h0007;
m[13'd5139]=16'h0000;
m[13'd5140]=16'h000e;
m[13'd5141]=16'h8104;
m[13'd5142]=16'h0060;
m[13'd5143]=16'h0003;
m[13'd5144]=16'h0009;
m[13'd5145]=16'h6002;
m[13'd5146]=16'h4bed;
m[13'd5147]=16'h000a;
m[13'd5148]=16'h0009;
m[13'd5149]=16'h7009;
m[13'd5150]=16'h0073;
m[13'd5151]=16'h0301;
m[13'd5152]=16'h0009;
m[13'd5153]=16'h9b00;
m[13'd5154]=16'h0018;
m[13'd5155]=16'h4104;
m[13'd5156]=16'h0060;
m[13'd5157]=16'h0003;
m[13'd5158]=16'h0009;
m[13'd5159]=16'h7002;
m[13'd5160]=16'h4bc0;
m[13'd5161]=16'h000a;
m[13'd5162]=16'h0009;
m[13'd5163]=16'h8009;
m[13'd5164]=16'h0073;
m[13'd5165]=16'h0301;
m[13'd5166]=16'h0009;
m[13'd5167]=16'h9b00;
m[13'd5168]=16'h0018;
m[13'd5169]=16'h4104;
m[13'd5170]=16'h0060;
m[13'd5171]=16'h0003;
m[13'd5172]=16'h0009;
m[13'd5173]=16'h8002;
m[13'd5174]=16'h4bc3;
m[13'd5175]=16'h000a;
m[13'd5176]=16'h0009;
m[13'd5177]=16'h9009;
m[13'd5178]=16'h0073;
m[13'd5179]=16'h0301;
m[13'd5180]=16'h0009;
m[13'd5181]=16'h9b00;
m[13'd5182]=16'h0018;
m[13'd5183]=16'h4104;
m[13'd5184]=16'h0060;
m[13'd5185]=16'h0003;
m[13'd5186]=16'h0009;
m[13'd5187]=16'h9002;
m[13'd5188]=16'h4bc3;
m[13'd5189]=16'h000a;
m[13'd5190]=16'h0009;
m[13'd5191]=16'ha009;
m[13'd5192]=16'h0073;
m[13'd5193]=16'h0301;
m[13'd5194]=16'h0009;
m[13'd5195]=16'h9b00;
m[13'd5196]=16'h0018;
m[13'd5197]=16'h4104;
m[13'd5198]=16'h0060;
m[13'd5199]=16'h0003;
m[13'd5200]=16'h0009;
m[13'd5201]=16'ha002;
m[13'd5202]=16'h4b95;
m[13'd5203]=16'h400b;
m[13'd5204]=16'h004e;
m[13'd5205]=16'h000a;
m[13'd5206]=16'h0009;
m[13'd5207]=16'hb009;
m[13'd5208]=16'h007b;
m[13'd5209]=16'h0301;
m[13'd5210]=16'h0009;
m[13'd5211]=16'h9b00;
m[13'd5212]=16'h0018;
m[13'd5213]=16'h4104;
m[13'd5214]=16'h0025;
m[13'd5215]=16'h4004;
m[13'd5216]=16'h004e;
m[13'd5217]=16'h0003;
m[13'd5218]=16'h0009;
m[13'd5219]=16'hb002;
m[13'd5220]=16'h4b4a;
m[13'd5221]=16'h400b;
m[13'd5222]=16'h004e;
m[13'd5223]=16'h000a;
m[13'd5224]=16'h0009;
m[13'd5225]=16'hc009;
m[13'd5226]=16'h0073;
m[13'd5227]=16'h0301;
m[13'd5228]=16'h0009;
m[13'd5229]=16'h9b00;
m[13'd5230]=16'h0018;
m[13'd5231]=16'h4104;
m[13'd5232]=16'h0025;
m[13'd5233]=16'h4004;
m[13'd5234]=16'h004e;
m[13'd5235]=16'h0003;
m[13'd5236]=16'h0009;
m[13'd5237]=16'hc002;
m[13'd5238]=16'h4b61;
m[13'd5239]=16'h400b;
m[13'd5240]=16'h004e;
m[13'd5241]=16'h000a;
m[13'd5242]=16'h0009;
m[13'd5243]=16'hd009;
m[13'd5244]=16'h0073;
m[13'd5245]=16'h0301;
m[13'd5246]=16'h0009;
m[13'd5247]=16'h9b00;
m[13'd5248]=16'h0018;
m[13'd5249]=16'h4104;
m[13'd5250]=16'h0025;
m[13'd5251]=16'h4004;
m[13'd5252]=16'h004e;
m[13'd5253]=16'h0003;
m[13'd5254]=16'h0009;
m[13'd5255]=16'hd002;
m[13'd5256]=16'h4b61;
m[13'd5257]=16'h400b;
m[13'd5258]=16'h004e;
m[13'd5259]=16'h000a;
m[13'd5260]=16'h0009;
m[13'd5261]=16'he009;
m[13'd5262]=16'h0073;
m[13'd5263]=16'h0301;
m[13'd5264]=16'h0009;
m[13'd5265]=16'h9b00;
m[13'd5266]=16'h0018;
m[13'd5267]=16'h4104;
m[13'd5268]=16'h0025;
m[13'd5269]=16'h4004;
m[13'd5270]=16'h004e;
m[13'd5271]=16'h0003;
m[13'd5272]=16'h0009;
m[13'd5273]=16'he002;
m[13'd5274]=16'h4b61;
m[13'd5275]=16'h400b;
m[13'd5276]=16'h004e;
m[13'd5277]=16'h000a;
m[13'd5278]=16'h0009;
m[13'd5279]=16'hf009;
m[13'd5280]=16'h0073;
m[13'd5281]=16'h0301;
m[13'd5282]=16'h0009;
m[13'd5283]=16'h9b00;
m[13'd5284]=16'h0018;
m[13'd5285]=16'h4104;
m[13'd5286]=16'h0025;
m[13'd5287]=16'h4004;
m[13'd5288]=16'h004e;
m[13'd5289]=16'h0003;
m[13'd5290]=16'h0009;
m[13'd5291]=16'hf002;
m[13'd5292]=16'h4b61;
m[13'd5293]=16'h400b;
m[13'd5294]=16'h004e;
m[13'd5295]=16'h010a;
m[13'd5296]=16'h0009;
m[13'd5297]=16'h0009;
m[13'd5298]=16'h0073;
m[13'd5299]=16'h0301;
m[13'd5300]=16'h0009;
m[13'd5301]=16'h9b00;
m[13'd5302]=16'h0018;
m[13'd5303]=16'h4104;
m[13'd5304]=16'h0025;
m[13'd5305]=16'h4004;
m[13'd5306]=16'h004e;
m[13'd5307]=16'h0103;
m[13'd5308]=16'h0009;
m[13'd5309]=16'h0002;
m[13'd5310]=16'h4be3;
m[13'd5311]=16'h0908;
m[13'd5312]=16'h0009;
m[13'd5313]=16'h9f07;
m[13'd5314]=16'h001b;
m[13'd5315]=16'h4009;
m[13'd5316]=16'h0010;
m[13'd5317]=16'h000a;
m[13'd5318]=16'h0016;
m[13'd5319]=16'h090c;
m[13'd5320]=16'h000a;
m[13'd5321]=16'h090d;
m[13'd5322]=16'h0007;
m[13'd5323]=16'h000b;
m[13'd5324]=16'h000a;
m[13'd5325]=16'h410b;
m[13'd5326]=16'h0095;
m[13'd5327]=16'h000a;
m[13'd5328]=16'h0009;
m[13'd5329]=16'h5009;
m[13'd5330]=16'h010f;
m[13'd5331]=16'h0301;
m[13'd5332]=16'h0009;
m[13'd5333]=16'h9b00;
m[13'd5334]=16'h001b;
m[13'd5335]=16'h4002;
m[13'd5336]=16'h0010;
m[13'd5337]=16'h0003;
m[13'd5338]=16'h0016;
m[13'd5339]=16'h0905;
m[13'd5340]=16'h000a;
m[13'd5341]=16'h0906;
m[13'd5342]=16'h0007;
m[13'd5343]=16'h0004;
m[13'd5344]=16'h000a;
m[13'd5345]=16'h4104;
m[13'd5346]=16'h008d;
m[13'd5347]=16'h0003;
m[13'd5348]=16'h0009;
m[13'd5349]=16'h5002;
m[13'd5350]=16'h4975;
m[13'd5351]=16'h000a;
m[13'd5352]=16'h0009;
m[13'd5353]=16'h6009;
m[13'd5354]=16'h0055;
m[13'd5355]=16'h4801;
m[13'd5356]=16'h0007;
m[13'd5357]=16'h0000;
m[13'd5358]=16'h000e;
m[13'd5359]=16'h8104;
m[13'd5360]=16'h0058;
m[13'd5361]=16'h0003;
m[13'd5362]=16'h0009;
m[13'd5363]=16'h6002;
m[13'd5364]=16'h4bf3;
m[13'd5365]=16'h000a;
m[13'd5366]=16'h0009;
m[13'd5367]=16'h7009;
m[13'd5368]=16'h0073;
m[13'd5369]=16'h0301;
m[13'd5370]=16'h0009;
m[13'd5371]=16'h9b00;
m[13'd5372]=16'h0018;
m[13'd5373]=16'h4104;
m[13'd5374]=16'h0058;
m[13'd5375]=16'h0003;
m[13'd5376]=16'h0009;
m[13'd5377]=16'h7002;
m[13'd5378]=16'h4bc9;
m[13'd5379]=16'h000a;
m[13'd5380]=16'h0009;
m[13'd5381]=16'h8009;
m[13'd5382]=16'h0073;
m[13'd5383]=16'h0301;
m[13'd5384]=16'h0009;
m[13'd5385]=16'h9b00;
m[13'd5386]=16'h0018;
m[13'd5387]=16'h4104;
m[13'd5388]=16'h0058;
m[13'd5389]=16'h0003;
m[13'd5390]=16'h0009;
m[13'd5391]=16'h8002;
m[13'd5392]=16'h4bcc;
m[13'd5393]=16'h000a;
m[13'd5394]=16'h0009;
m[13'd5395]=16'h9009;
m[13'd5396]=16'h0073;
m[13'd5397]=16'h0301;
m[13'd5398]=16'h0009;
m[13'd5399]=16'h9b00;
m[13'd5400]=16'h0018;
m[13'd5401]=16'h4104;
m[13'd5402]=16'h0058;
m[13'd5403]=16'h0003;
m[13'd5404]=16'h0009;
m[13'd5405]=16'h9002;
m[13'd5406]=16'h4bc9;
m[13'd5407]=16'h000a;
m[13'd5408]=16'h0009;
m[13'd5409]=16'ha009;
m[13'd5410]=16'h0073;
m[13'd5411]=16'h0301;
m[13'd5412]=16'h0009;
m[13'd5413]=16'h9b00;
m[13'd5414]=16'h0018;
m[13'd5415]=16'h4104;
m[13'd5416]=16'h0058;
m[13'd5417]=16'h0003;
m[13'd5418]=16'h0009;
m[13'd5419]=16'ha002;
m[13'd5420]=16'h4b9e;
m[13'd5421]=16'h400b;
m[13'd5422]=16'h004e;
m[13'd5423]=16'h000a;
m[13'd5424]=16'h0009;
m[13'd5425]=16'hb009;
m[13'd5426]=16'h0102;
m[13'd5427]=16'h0401;
m[13'd5428]=16'h0009;
m[13'd5429]=16'hd000;
m[13'd5430]=16'h001b;
m[13'd5431]=16'h4002;
m[13'd5432]=16'h0010;
m[13'd5433]=16'h0003;
m[13'd5434]=16'h0016;
m[13'd5435]=16'h0905;
m[13'd5436]=16'h000a;
m[13'd5437]=16'h0906;
m[13'd5438]=16'h0007;
m[13'd5439]=16'h0004;
m[13'd5440]=16'h000a;
m[13'd5441]=16'h4104;
m[13'd5442]=16'h008d;
m[13'd5443]=16'h0003;
m[13'd5444]=16'h0009;
m[13'd5445]=16'h5002;
m[13'd5446]=16'h4a66;
m[13'd5447]=16'h400b;
m[13'd5448]=16'h004e;
m[13'd5449]=16'h000a;
m[13'd5450]=16'h0009;
m[13'd5451]=16'hc009;
m[13'd5452]=16'h0055;
m[13'd5453]=16'h4801;
m[13'd5454]=16'h0007;
m[13'd5455]=16'h0000;
m[13'd5456]=16'h000e;
m[13'd5457]=16'h8104;
m[13'd5458]=16'h0058;
m[13'd5459]=16'h0003;
m[13'd5460]=16'h0009;
m[13'd5461]=16'h6002;
m[13'd5462]=16'h4ba6;
m[13'd5463]=16'h400b;
m[13'd5464]=16'h004e;
m[13'd5465]=16'h000a;
m[13'd5466]=16'h0009;
m[13'd5467]=16'hd009;
m[13'd5468]=16'h0073;
m[13'd5469]=16'h0401;
m[13'd5470]=16'h0009;
m[13'd5471]=16'hd000;
m[13'd5472]=16'h0018;
m[13'd5473]=16'h4104;
m[13'd5474]=16'h0058;
m[13'd5475]=16'h0003;
m[13'd5476]=16'h0009;
m[13'd5477]=16'h7002;
m[13'd5478]=16'h4b7c;
m[13'd5479]=16'h400b;
m[13'd5480]=16'h004e;
m[13'd5481]=16'h000a;
m[13'd5482]=16'h0009;
m[13'd5483]=16'he009;
m[13'd5484]=16'h0073;
m[13'd5485]=16'h0401;
m[13'd5486]=16'h0009;
m[13'd5487]=16'hd000;
m[13'd5488]=16'h0018;
m[13'd5489]=16'h4104;
m[13'd5490]=16'h0058;
m[13'd5491]=16'h0003;
m[13'd5492]=16'h0009;
m[13'd5493]=16'h8002;
m[13'd5494]=16'h4b7c;
m[13'd5495]=16'h400b;
m[13'd5496]=16'h004e;
m[13'd5497]=16'h000a;
m[13'd5498]=16'h0009;
m[13'd5499]=16'hf009;
m[13'd5500]=16'h0073;
m[13'd5501]=16'h0401;
m[13'd5502]=16'h0009;
m[13'd5503]=16'hd000;
m[13'd5504]=16'h0018;
m[13'd5505]=16'h4104;
m[13'd5506]=16'h0058;
m[13'd5507]=16'h0003;
m[13'd5508]=16'h0009;
m[13'd5509]=16'h9002;
m[13'd5510]=16'h4b7c;
m[13'd5511]=16'h400b;
m[13'd5512]=16'h004e;
m[13'd5513]=16'h010a;
m[13'd5514]=16'h0009;
m[13'd5515]=16'h0009;
m[13'd5516]=16'h0073;
m[13'd5517]=16'h0401;
m[13'd5518]=16'h0009;
m[13'd5519]=16'hd000;
m[13'd5520]=16'h0018;
m[13'd5521]=16'h4104;
m[13'd5522]=16'h0058;
m[13'd5523]=16'h0003;
m[13'd5524]=16'h0009;
m[13'd5525]=16'ha002;
m[13'd5526]=16'h4bc7;
m[13'd5527]=16'h010a;
m[13'd5528]=16'h0009;
m[13'd5529]=16'h1009;
m[13'd5530]=16'h0102;
m[13'd5531]=16'h0301;
m[13'd5532]=16'h0009;
m[13'd5533]=16'h9b00;
m[13'd5534]=16'h001b;
m[13'd5535]=16'h4002;
m[13'd5536]=16'h0010;
m[13'd5537]=16'h0003;
m[13'd5538]=16'h0016;
m[13'd5539]=16'h0905;
m[13'd5540]=16'h000a;
m[13'd5541]=16'h0906;
m[13'd5542]=16'h0007;
m[13'd5543]=16'h0004;
m[13'd5544]=16'h000a;
m[13'd5545]=16'h4104;
m[13'd5546]=16'h008d;
m[13'd5547]=16'h0003;
m[13'd5548]=16'h0009;
m[13'd5549]=16'h5002;
m[13'd5550]=16'h4ab0;
m[13'd5551]=16'h010a;
m[13'd5552]=16'h0009;
m[13'd5553]=16'h2009;
m[13'd5554]=16'h0055;
m[13'd5555]=16'h4801;
m[13'd5556]=16'h0007;
m[13'd5557]=16'h0000;
m[13'd5558]=16'h000e;
m[13'd5559]=16'h8104;
m[13'd5560]=16'h0058;
m[13'd5561]=16'h0003;
m[13'd5562]=16'h0009;
m[13'd5563]=16'h6002;
m[13'd5564]=16'h4bf6;
m[13'd5565]=16'h010a;
m[13'd5566]=16'h0009;
m[13'd5567]=16'h3009;
m[13'd5568]=16'h0073;
m[13'd5569]=16'h0301;
m[13'd5570]=16'h0009;
m[13'd5571]=16'h9b00;
m[13'd5572]=16'h0018;
m[13'd5573]=16'h4104;
m[13'd5574]=16'h0058;
m[13'd5575]=16'h0003;
m[13'd5576]=16'h0009;
m[13'd5577]=16'h7002;
m[13'd5578]=16'h4bc9;
m[13'd5579]=16'h010a;
m[13'd5580]=16'h0009;
m[13'd5581]=16'h4009;
m[13'd5582]=16'h0073;
m[13'd5583]=16'h0301;
m[13'd5584]=16'h0009;
m[13'd5585]=16'h9b00;
m[13'd5586]=16'h0018;
m[13'd5587]=16'h4104;
m[13'd5588]=16'h0058;
m[13'd5589]=16'h0003;
m[13'd5590]=16'h0009;
m[13'd5591]=16'h8002;
m[13'd5592]=16'h4bc9;
m[13'd5593]=16'h010a;
m[13'd5594]=16'h0009;
m[13'd5595]=16'h5009;
m[13'd5596]=16'h0073;
m[13'd5597]=16'h0301;
m[13'd5598]=16'h0009;
m[13'd5599]=16'h9b00;
m[13'd5600]=16'h0018;
m[13'd5601]=16'h4104;
m[13'd5602]=16'h0058;
m[13'd5603]=16'h0003;
m[13'd5604]=16'h0009;
m[13'd5605]=16'h9002;
m[13'd5606]=16'h4bcc;
m[13'd5607]=16'h010a;
m[13'd5608]=16'h0009;
m[13'd5609]=16'h6009;
m[13'd5610]=16'h0073;
m[13'd5611]=16'h0301;
m[13'd5612]=16'h0009;
m[13'd5613]=16'h9b00;
m[13'd5614]=16'h0018;
m[13'd5615]=16'h4104;
m[13'd5616]=16'h0058;
m[13'd5617]=16'h0003;
m[13'd5618]=16'h0009;
m[13'd5619]=16'ha002;
m[13'd5620]=16'h4c10;
m[13'd5621]=16'h0808;
m[13'd5622]=16'h0009;
m[13'd5623]=16'h9307;
m[13'd5624]=16'h001b;
m[13'd5625]=16'h4009;
m[13'd5626]=16'h0010;
m[13'd5627]=16'h000a;
m[13'd5628]=16'h0016;
m[13'd5629]=16'h090c;
m[13'd5630]=16'h000a;
m[13'd5631]=16'h090d;
m[13'd5632]=16'h0007;
m[13'd5633]=16'h000b;
m[13'd5634]=16'h000a;
m[13'd5635]=16'h410b;
m[13'd5636]=16'h008d;
m[13'd5637]=16'h000a;
m[13'd5638]=16'h0009;
m[13'd5639]=16'h5009;
m[13'd5640]=16'h0102;
m[13'd5641]=16'h0301;
m[13'd5642]=16'h0009;
m[13'd5643]=16'h9b00;
m[13'd5644]=16'h001b;
m[13'd5645]=16'h4002;
m[13'd5646]=16'h0010;
m[13'd5647]=16'h0003;
m[13'd5648]=16'h0016;
m[13'd5649]=16'h0905;
m[13'd5650]=16'h000a;
m[13'd5651]=16'h0906;
m[13'd5652]=16'h0007;
m[13'd5653]=16'h0004;
m[13'd5654]=16'h000a;
m[13'd5655]=16'h4104;
m[13'd5656]=16'h008d;
m[13'd5657]=16'h0003;
m[13'd5658]=16'h0009;
m[13'd5659]=16'h5002;
m[13'd5660]=16'h4982;
m[13'd5661]=16'h000a;
m[13'd5662]=16'h0009;
m[13'd5663]=16'h6009;
m[13'd5664]=16'h0055;
m[13'd5665]=16'h4801;
m[13'd5666]=16'h0007;
m[13'd5667]=16'h0000;
m[13'd5668]=16'h000e;
m[13'd5669]=16'h8104;
m[13'd5670]=16'h0058;
m[13'd5671]=16'h0003;
m[13'd5672]=16'h0009;
m[13'd5673]=16'h6002;
m[13'd5674]=16'h4bf4;
m[13'd5675]=16'h000a;
m[13'd5676]=16'h0009;
m[13'd5677]=16'h7009;
m[13'd5678]=16'h0073;
m[13'd5679]=16'h0301;
m[13'd5680]=16'h0009;
m[13'd5681]=16'h9b00;
m[13'd5682]=16'h0018;
m[13'd5683]=16'h4104;
m[13'd5684]=16'h0058;
m[13'd5685]=16'h0003;
m[13'd5686]=16'h0009;
m[13'd5687]=16'h7002;
m[13'd5688]=16'h4bca;
m[13'd5689]=16'h000a;
m[13'd5690]=16'h0009;
m[13'd5691]=16'h8009;
m[13'd5692]=16'h0073;
m[13'd5693]=16'h0301;
m[13'd5694]=16'h0009;
m[13'd5695]=16'h9b00;
m[13'd5696]=16'h0018;
m[13'd5697]=16'h4104;
m[13'd5698]=16'h0058;
m[13'd5699]=16'h0003;
m[13'd5700]=16'h0009;
m[13'd5701]=16'h8002;
m[13'd5702]=16'h4bca;
m[13'd5703]=16'h000a;
m[13'd5704]=16'h0009;
m[13'd5705]=16'h9009;
m[13'd5706]=16'h0073;
m[13'd5707]=16'h0301;
m[13'd5708]=16'h0009;
m[13'd5709]=16'h9b00;
m[13'd5710]=16'h0018;
m[13'd5711]=16'h4104;
m[13'd5712]=16'h0058;
m[13'd5713]=16'h0003;
m[13'd5714]=16'h0009;
m[13'd5715]=16'h9002;
m[13'd5716]=16'h4bca;
m[13'd5717]=16'h000a;
m[13'd5718]=16'h0009;
m[13'd5719]=16'ha009;
m[13'd5720]=16'h0073;
m[13'd5721]=16'h0301;
m[13'd5722]=16'h0009;
m[13'd5723]=16'h9b00;
m[13'd5724]=16'h0018;
m[13'd5725]=16'h4104;
m[13'd5726]=16'h0058;
m[13'd5727]=16'h0003;
m[13'd5728]=16'h0009;
m[13'd5729]=16'ha002;
m[13'd5730]=16'h4c2f;
m[13'd5731]=16'h0108;
m[13'd5732]=16'h0009;
m[13'd5733]=16'h2307;
m[13'd5734]=16'h001b;
m[13'd5735]=16'h4009;
m[13'd5736]=16'h0010;
m[13'd5737]=16'h000a;
m[13'd5738]=16'h0016;
m[13'd5739]=16'h090c;
m[13'd5740]=16'h000a;
m[13'd5741]=16'h090d;
m[13'd5742]=16'h0007;
m[13'd5743]=16'h000b;
m[13'd5744]=16'h000a;
m[13'd5745]=16'h410b;
m[13'd5746]=16'h0095;
m[13'd5747]=16'h000a;
m[13'd5748]=16'h0009;
m[13'd5749]=16'h5009;
m[13'd5750]=16'h0102;
m[13'd5751]=16'h0401;
m[13'd5752]=16'h0009;
m[13'd5753]=16'h4900;
m[13'd5754]=16'h001b;
m[13'd5755]=16'h4002;
m[13'd5756]=16'h0010;
m[13'd5757]=16'h0003;
m[13'd5758]=16'h0016;
m[13'd5759]=16'h0905;
m[13'd5760]=16'h000a;
m[13'd5761]=16'h0906;
m[13'd5762]=16'h0007;
m[13'd5763]=16'h0004;
m[13'd5764]=16'h000a;
m[13'd5765]=16'h4104;
m[13'd5766]=16'h008d;
m[13'd5767]=16'h0003;
m[13'd5768]=16'h0009;
m[13'd5769]=16'h5002;
m[13'd5770]=16'h4930;
m[13'd5771]=16'h810b;
m[13'd5772]=16'h002b;
m[13'd5773]=16'h3108;
m[13'd5774]=16'h0007;
m[13'd5775]=16'h0007;
m[13'd5776]=16'h0060;
m[13'd5777]=16'h000a;
m[13'd5778]=16'h0009;
m[13'd5779]=16'h6009;
m[13'd5780]=16'h0055;
m[13'd5781]=16'h4801;
m[13'd5782]=16'h0007;
m[13'd5783]=16'h0000;
m[13'd5784]=16'h000e;
m[13'd5785]=16'h8104;
m[13'd5786]=16'h0058;
m[13'd5787]=16'h0003;
m[13'd5788]=16'h0009;
m[13'd5789]=16'h6002;
m[13'd5790]=16'h4b63;
m[13'd5791]=16'h110b;
m[13'd5792]=16'h002b;
m[13'd5793]=16'h1108;
m[13'd5794]=16'h0007;
m[13'd5795]=16'h0007;
m[13'd5796]=16'h0060;
m[13'd5797]=16'h000a;
m[13'd5798]=16'h0009;
m[13'd5799]=16'h7009;
m[13'd5800]=16'h0073;
m[13'd5801]=16'h0401;
m[13'd5802]=16'h0009;
m[13'd5803]=16'h4900;
m[13'd5804]=16'h0018;
m[13'd5805]=16'h4104;
m[13'd5806]=16'h0058;
m[13'd5807]=16'h0003;
m[13'd5808]=16'h0009;
m[13'd5809]=16'h7002;
m[13'd5810]=16'h4b39;
m[13'd5811]=16'h800b;
m[13'd5812]=16'h002b;
m[13'd5813]=16'h0808;
m[13'd5814]=16'h0007;
m[13'd5815]=16'h0007;
m[13'd5816]=16'h0060;
m[13'd5817]=16'h000a;
m[13'd5818]=16'h0009;
m[13'd5819]=16'h8009;
m[13'd5820]=16'h0073;
m[13'd5821]=16'h0401;
m[13'd5822]=16'h0009;
m[13'd5823]=16'h4900;
m[13'd5824]=16'h0018;
m[13'd5825]=16'h4104;
m[13'd5826]=16'h0058;
m[13'd5827]=16'h0003;
m[13'd5828]=16'h0009;
m[13'd5829]=16'h8002;
m[13'd5830]=16'h4b36;
m[13'd5831]=16'h400b;
m[13'd5832]=16'h002b;
m[13'd5833]=16'h1608;
m[13'd5834]=16'h0007;
m[13'd5835]=16'h0007;
m[13'd5836]=16'h0060;
m[13'd5837]=16'h000a;
m[13'd5838]=16'h0009;
m[13'd5839]=16'h9009;
m[13'd5840]=16'h0073;
m[13'd5841]=16'h0401;
m[13'd5842]=16'h0009;
m[13'd5843]=16'h4900;
m[13'd5844]=16'h0018;
m[13'd5845]=16'h4104;
m[13'd5846]=16'h0058;
m[13'd5847]=16'h0003;
m[13'd5848]=16'h0009;
m[13'd5849]=16'h9002;
m[13'd5850]=16'h4b39;
m[13'd5851]=16'h800b;
m[13'd5852]=16'h002b;
m[13'd5853]=16'h0508;
m[13'd5854]=16'h0007;
m[13'd5855]=16'h0007;
m[13'd5856]=16'h0060;
m[13'd5857]=16'h000a;
m[13'd5858]=16'h0009;
m[13'd5859]=16'ha009;
m[13'd5860]=16'h0073;
m[13'd5861]=16'h0401;
m[13'd5862]=16'h0009;
m[13'd5863]=16'h4900;
m[13'd5864]=16'h0018;
m[13'd5865]=16'h4104;
m[13'd5866]=16'h0058;
m[13'd5867]=16'h0003;
m[13'd5868]=16'h0009;
m[13'd5869]=16'ha002;
m[13'd5870]=16'h4b49;
m[13'd5871]=16'h800b;
m[13'd5872]=16'h002b;
m[13'd5873]=16'h0408;
m[13'd5874]=16'h0007;
m[13'd5875]=16'h0007;
m[13'd5876]=16'h0025;
m[13'd5877]=16'h400b;
m[13'd5878]=16'h004e;
m[13'd5879]=16'h000a;
m[13'd5880]=16'h0009;
m[13'd5881]=16'hb009;
m[13'd5882]=16'h010f;
m[13'd5883]=16'h0301;
m[13'd5884]=16'h0009;
m[13'd5885]=16'h9b00;
m[13'd5886]=16'h001b;
m[13'd5887]=16'h4002;
m[13'd5888]=16'h0010;
m[13'd5889]=16'h0003;
m[13'd5890]=16'h0016;
m[13'd5891]=16'h0905;
m[13'd5892]=16'h000a;
m[13'd5893]=16'h0906;
m[13'd5894]=16'h0007;
m[13'd5895]=16'h0004;
m[13'd5896]=16'h000a;
m[13'd5897]=16'h4104;
m[13'd5898]=16'h0095;
m[13'd5899]=16'h0003;
m[13'd5900]=16'h0009;
m[13'd5901]=16'h5002;
m[13'd5902]=16'h49f6;
m[13'd5903]=16'h800b;
m[13'd5904]=16'h002b;
m[13'd5905]=16'h0308;
m[13'd5906]=16'h0007;
m[13'd5907]=16'h0007;
m[13'd5908]=16'h0025;
m[13'd5909]=16'h400b;
m[13'd5910]=16'h004e;
m[13'd5911]=16'h000a;
m[13'd5912]=16'h0009;
m[13'd5913]=16'hc009;
m[13'd5914]=16'h0055;
m[13'd5915]=16'h4801;
m[13'd5916]=16'h0007;
m[13'd5917]=16'h0000;
m[13'd5918]=16'h000e;
m[13'd5919]=16'h8104;
m[13'd5920]=16'h0060;
m[13'd5921]=16'h0003;
m[13'd5922]=16'h0009;
m[13'd5923]=16'h6002;
m[13'd5924]=16'h4b48;
m[13'd5925]=16'h800b;
m[13'd5926]=16'h002b;
m[13'd5927]=16'h0308;
m[13'd5928]=16'h0007;
m[13'd5929]=16'h0007;
m[13'd5930]=16'h0025;
m[13'd5931]=16'h400b;
m[13'd5932]=16'h004e;
m[13'd5933]=16'h000a;
m[13'd5934]=16'h0009;
m[13'd5935]=16'hd009;
m[13'd5936]=16'h0073;
m[13'd5937]=16'h0301;
m[13'd5938]=16'h0009;
m[13'd5939]=16'h9b00;
m[13'd5940]=16'h0018;
m[13'd5941]=16'h4104;
m[13'd5942]=16'h0060;
m[13'd5943]=16'h0003;
m[13'd5944]=16'h0009;
m[13'd5945]=16'h7002;
m[13'd5946]=16'h4b1e;
m[13'd5947]=16'h100b;
m[13'd5948]=16'h002b;
m[13'd5949]=16'h1208;
m[13'd5950]=16'h0007;
m[13'd5951]=16'h0007;
m[13'd5952]=16'h0025;
m[13'd5953]=16'h400b;
m[13'd5954]=16'h004e;
m[13'd5955]=16'h000a;
m[13'd5956]=16'h0009;
m[13'd5957]=16'he009;
m[13'd5958]=16'h0073;
m[13'd5959]=16'h0301;
m[13'd5960]=16'h0009;
m[13'd5961]=16'h9b00;
m[13'd5962]=16'h0018;
m[13'd5963]=16'h4104;
m[13'd5964]=16'h0060;
m[13'd5965]=16'h0003;
m[13'd5966]=16'h0009;
m[13'd5967]=16'h8002;
m[13'd5968]=16'h4b1b;
m[13'd5969]=16'h100b;
m[13'd5970]=16'h002b;
m[13'd5971]=16'h1208;
m[13'd5972]=16'h0007;
m[13'd5973]=16'h0007;
m[13'd5974]=16'h0025;
m[13'd5975]=16'h400b;
m[13'd5976]=16'h004e;
m[13'd5977]=16'h000a;
m[13'd5978]=16'h0009;
m[13'd5979]=16'hf009;
m[13'd5980]=16'h0073;
m[13'd5981]=16'h0301;
m[13'd5982]=16'h0009;
m[13'd5983]=16'h9b00;
m[13'd5984]=16'h0018;
m[13'd5985]=16'h4104;
m[13'd5986]=16'h0060;
m[13'd5987]=16'h0003;
m[13'd5988]=16'h0009;
m[13'd5989]=16'h9002;
m[13'd5990]=16'h4b1e;
m[13'd5991]=16'h100b;
m[13'd5992]=16'h002b;
m[13'd5993]=16'h1108;
m[13'd5994]=16'h0007;
m[13'd5995]=16'h0007;
m[13'd5996]=16'h0025;
m[13'd5997]=16'h400b;
m[13'd5998]=16'h004e;
m[13'd5999]=16'h010a;
m[13'd6000]=16'h0009;
m[13'd6001]=16'h0009;
m[13'd6002]=16'h0073;
m[13'd6003]=16'h0301;
m[13'd6004]=16'h0009;
m[13'd6005]=16'h9b00;
m[13'd6006]=16'h0018;
m[13'd6007]=16'h4104;
m[13'd6008]=16'h0060;
m[13'd6009]=16'h0003;
m[13'd6010]=16'h0009;
m[13'd6011]=16'ha002;
m[13'd6012]=16'h4ba8;
m[13'd6013]=16'h0608;
m[13'd6014]=16'h0009;
m[13'd6015]=16'h6c07;
m[13'd6016]=16'h001b;
m[13'd6017]=16'h4009;
m[13'd6018]=16'h0010;
m[13'd6019]=16'h000a;
m[13'd6020]=16'h0016;
m[13'd6021]=16'h090c;
m[13'd6022]=16'h000a;
m[13'd6023]=16'h090d;
m[13'd6024]=16'h0007;
m[13'd6025]=16'h000b;
m[13'd6026]=16'h000a;
m[13'd6027]=16'h410b;
m[13'd6028]=16'h0095;
m[13'd6029]=16'h000a;
m[13'd6030]=16'h0009;
m[13'd6031]=16'h5009;
m[13'd6032]=16'h007b;
m[13'd6033]=16'h0301;
m[13'd6034]=16'h0009;
m[13'd6035]=16'h9b00;
m[13'd6036]=16'h0018;
m[13'd6037]=16'h4104;
m[13'd6038]=16'h0025;
m[13'd6039]=16'h4004;
m[13'd6040]=16'h004e;
m[13'd6041]=16'h0003;
m[13'd6042]=16'h0009;
m[13'd6043]=16'hb002;
m[13'd6044]=16'h4a5c;
m[13'd6045]=16'h000a;
m[13'd6046]=16'h0009;
m[13'd6047]=16'h6009;
m[13'd6048]=16'h0073;
m[13'd6049]=16'h0301;
m[13'd6050]=16'h0009;
m[13'd6051]=16'h9b00;
m[13'd6052]=16'h0018;
m[13'd6053]=16'h4104;
m[13'd6054]=16'h0025;
m[13'd6055]=16'h4004;
m[13'd6056]=16'h004e;
m[13'd6057]=16'h0003;
m[13'd6058]=16'h0009;
m[13'd6059]=16'hc002;
m[13'd6060]=16'h4bae;
m[13'd6061]=16'h000a;
m[13'd6062]=16'h0009;
m[13'd6063]=16'h7009;
m[13'd6064]=16'h0073;
m[13'd6065]=16'h0301;
m[13'd6066]=16'h0009;
m[13'd6067]=16'h9b00;
m[13'd6068]=16'h0018;
m[13'd6069]=16'h4104;
m[13'd6070]=16'h0025;
m[13'd6071]=16'h4004;
m[13'd6072]=16'h004e;
m[13'd6073]=16'h0003;
m[13'd6074]=16'h0009;
m[13'd6075]=16'hd002;
m[13'd6076]=16'h4bae;
m[13'd6077]=16'h000a;
m[13'd6078]=16'h0009;
m[13'd6079]=16'h8009;
m[13'd6080]=16'h0073;
m[13'd6081]=16'h0301;
m[13'd6082]=16'h0009;
m[13'd6083]=16'h9b00;
m[13'd6084]=16'h0018;
m[13'd6085]=16'h4104;
m[13'd6086]=16'h0025;
m[13'd6087]=16'h4004;
m[13'd6088]=16'h004e;
m[13'd6089]=16'h0003;
m[13'd6090]=16'h0009;
m[13'd6091]=16'he002;
m[13'd6092]=16'h4bb1;
m[13'd6093]=16'h000a;
m[13'd6094]=16'h0009;
m[13'd6095]=16'h9009;
m[13'd6096]=16'h0073;
m[13'd6097]=16'h0301;
m[13'd6098]=16'h0009;
m[13'd6099]=16'h9b00;
m[13'd6100]=16'h0018;
m[13'd6101]=16'h4104;
m[13'd6102]=16'h0025;
m[13'd6103]=16'h4004;
m[13'd6104]=16'h004e;
m[13'd6105]=16'h0003;
m[13'd6106]=16'h0009;
m[13'd6107]=16'hf002;
m[13'd6108]=16'h4bae;
m[13'd6109]=16'h000a;
m[13'd6110]=16'h0009;
m[13'd6111]=16'ha009;
m[13'd6112]=16'h0073;
m[13'd6113]=16'h0301;
m[13'd6114]=16'h0009;
m[13'd6115]=16'h9b00;
m[13'd6116]=16'h0018;
m[13'd6117]=16'h4104;
m[13'd6118]=16'h0025;
m[13'd6119]=16'h4004;
m[13'd6120]=16'h004e;
m[13'd6121]=16'h0103;
m[13'd6122]=16'h0009;
m[13'd6123]=16'h0002;
m[13'd6124]=16'h4b83;
m[13'd6125]=16'h400b;
m[13'd6126]=16'h004e;
m[13'd6127]=16'h000a;
m[13'd6128]=16'h0009;
m[13'd6129]=16'hb009;
m[13'd6130]=16'h010f;
m[13'd6131]=16'h0301;
m[13'd6132]=16'h0009;
m[13'd6133]=16'h3600;
m[13'd6134]=16'h001b;
m[13'd6135]=16'h4002;
m[13'd6136]=16'h0010;
m[13'd6137]=16'h0003;
m[13'd6138]=16'h0016;
m[13'd6139]=16'h0905;
m[13'd6140]=16'h000a;
m[13'd6141]=16'h0906;
m[13'd6142]=16'h0007;
m[13'd6143]=16'h0004;
m[13'd6144]=16'h000a;
m[13'd6145]=16'h4104;
m[13'd6146]=16'h008d;
m[13'd6147]=16'h0003;
m[13'd6148]=16'h0009;
m[13'd6149]=16'h5002;
m[13'd6150]=16'h4a57;
m[13'd6151]=16'h400b;
m[13'd6152]=16'h004e;
m[13'd6153]=16'h000a;
m[13'd6154]=16'h0009;
m[13'd6155]=16'hc009;
m[13'd6156]=16'h0055;
m[13'd6157]=16'h4801;
m[13'd6158]=16'h0007;
m[13'd6159]=16'h0000;
m[13'd6160]=16'h000e;
m[13'd6161]=16'h8104;
m[13'd6162]=16'h0058;
m[13'd6163]=16'h0003;
m[13'd6164]=16'h0009;
m[13'd6165]=16'h6002;
m[13'd6166]=16'h4ba6;
m[13'd6167]=16'h400b;
m[13'd6168]=16'h004e;
m[13'd6169]=16'h000a;
m[13'd6170]=16'h0009;
m[13'd6171]=16'hd009;
m[13'd6172]=16'h0073;
m[13'd6173]=16'h0301;
m[13'd6174]=16'h0009;
m[13'd6175]=16'h3600;
m[13'd6176]=16'h0018;
m[13'd6177]=16'h4104;
m[13'd6178]=16'h0058;
m[13'd6179]=16'h0003;
m[13'd6180]=16'h0009;
m[13'd6181]=16'h7002;
m[13'd6182]=16'h4b7c;
m[13'd6183]=16'h400b;
m[13'd6184]=16'h004e;
m[13'd6185]=16'h000a;
m[13'd6186]=16'h0009;
m[13'd6187]=16'he009;
m[13'd6188]=16'h0073;
m[13'd6189]=16'h0301;
m[13'd6190]=16'h0009;
m[13'd6191]=16'h3600;
m[13'd6192]=16'h0018;
m[13'd6193]=16'h4104;
m[13'd6194]=16'h0058;
m[13'd6195]=16'h0003;
m[13'd6196]=16'h0009;
m[13'd6197]=16'h8002;
m[13'd6198]=16'h4b7c;
m[13'd6199]=16'h400b;
m[13'd6200]=16'h004e;
m[13'd6201]=16'h000a;
m[13'd6202]=16'h0009;
m[13'd6203]=16'hf009;
m[13'd6204]=16'h0073;
m[13'd6205]=16'h0301;
m[13'd6206]=16'h0009;
m[13'd6207]=16'h3600;
m[13'd6208]=16'h0018;
m[13'd6209]=16'h4104;
m[13'd6210]=16'h0058;
m[13'd6211]=16'h0003;
m[13'd6212]=16'h0009;
m[13'd6213]=16'h9002;
m[13'd6214]=16'h4b7c;
m[13'd6215]=16'h400b;
m[13'd6216]=16'h004e;
m[13'd6217]=16'h010a;
m[13'd6218]=16'h0009;
m[13'd6219]=16'h0009;
m[13'd6220]=16'h0073;
m[13'd6221]=16'h0301;
m[13'd6222]=16'h0009;
m[13'd6223]=16'h3600;
m[13'd6224]=16'h0018;
m[13'd6225]=16'h4104;
m[13'd6226]=16'h0058;
m[13'd6227]=16'h0003;
m[13'd6228]=16'h0009;
m[13'd6229]=16'ha002;
m[13'd6230]=16'h4af5;
m[13'd6231]=16'h4012;
m[13'd6232]=16'h0199;
m[13'd6233]=16'h0708;
m[13'd6234]=16'h0009;
m[13'd6235]=16'h3507;
m[13'd6236]=16'h001b;
m[13'd6237]=16'h4009;
m[13'd6238]=16'h0010;
m[13'd6239]=16'h000a;
m[13'd6240]=16'h0016;
m[13'd6241]=16'h090c;
m[13'd6242]=16'h000a;
m[13'd6243]=16'h090d;
m[13'd6244]=16'h0007;
m[13'd6245]=16'h000b;
m[13'd6246]=16'h000a;
m[13'd6247]=16'h410b;
m[13'd6248]=16'h0095;
m[13'd6249]=16'h000a;
m[13'd6250]=16'h0009;
m[13'd6251]=16'h5009;
m[13'd6252]=16'h010f;
m[13'd6253]=16'h0301;
m[13'd6254]=16'h0009;
m[13'd6255]=16'h9b00;
m[13'd6256]=16'h001b;
m[13'd6257]=16'h4002;
m[13'd6258]=16'h0010;
m[13'd6259]=16'h0003;
m[13'd6260]=16'h0016;
m[13'd6261]=16'h0905;
m[13'd6262]=16'h000a;
m[13'd6263]=16'h0906;
m[13'd6264]=16'h0007;
m[13'd6265]=16'h0004;
m[13'd6266]=16'h000a;
m[13'd6267]=16'h4104;
m[13'd6268]=16'h0095;
m[13'd6269]=16'h0003;
m[13'd6270]=16'h0009;
m[13'd6271]=16'h5002;
m[13'd6272]=16'h4812;
m[13'd6273]=16'h4012;
m[13'd6274]=16'h00dc;
m[13'd6275]=16'h000a;
m[13'd6276]=16'h0009;
m[13'd6277]=16'h6009;
m[13'd6278]=16'h0055;
m[13'd6279]=16'h4801;
m[13'd6280]=16'h0007;
m[13'd6281]=16'h0000;
m[13'd6282]=16'h000e;
m[13'd6283]=16'h8104;
m[13'd6284]=16'h0060;
m[13'd6285]=16'h0003;
m[13'd6286]=16'h0009;
m[13'd6287]=16'h6002;
m[13'd6288]=16'h4b11;
m[13'd6289]=16'h4012;
m[13'd6290]=16'h00dc;
m[13'd6291]=16'h000a;
m[13'd6292]=16'h0009;
m[13'd6293]=16'h7009;
m[13'd6294]=16'h0073;
m[13'd6295]=16'h0301;
m[13'd6296]=16'h0009;
m[13'd6297]=16'h9b00;
m[13'd6298]=16'h0018;
m[13'd6299]=16'h4104;
m[13'd6300]=16'h0060;
m[13'd6301]=16'h0003;
m[13'd6302]=16'h0009;
m[13'd6303]=16'h7002;
m[13'd6304]=16'h4ae7;
m[13'd6305]=16'h4012;
m[13'd6306]=16'h00dc;
m[13'd6307]=16'h000a;
m[13'd6308]=16'h0009;
m[13'd6309]=16'h8009;
m[13'd6310]=16'h0073;
m[13'd6311]=16'h0301;
m[13'd6312]=16'h0009;
m[13'd6313]=16'h9b00;
m[13'd6314]=16'h0018;
m[13'd6315]=16'h4104;
m[13'd6316]=16'h0060;
m[13'd6317]=16'h0003;
m[13'd6318]=16'h0009;
m[13'd6319]=16'h8002;
m[13'd6320]=16'h4ae4;
m[13'd6321]=16'h4012;
m[13'd6322]=16'h00dc;
m[13'd6323]=16'h000a;
m[13'd6324]=16'h0009;
m[13'd6325]=16'h9009;
m[13'd6326]=16'h0073;
m[13'd6327]=16'h0301;
m[13'd6328]=16'h0009;
m[13'd6329]=16'h9b00;
m[13'd6330]=16'h0018;
m[13'd6331]=16'h4104;
m[13'd6332]=16'h0060;
m[13'd6333]=16'h0003;
m[13'd6334]=16'h0009;
m[13'd6335]=16'h9002;
m[13'd6336]=16'h4ae7;
m[13'd6337]=16'h4012;
m[13'd6338]=16'h00dc;
m[13'd6339]=16'h000a;
m[13'd6340]=16'h0009;
m[13'd6341]=16'ha009;
m[13'd6342]=16'h0073;
m[13'd6343]=16'h0301;
m[13'd6344]=16'h0009;
m[13'd6345]=16'h9b00;
m[13'd6346]=16'h0018;
m[13'd6347]=16'h4104;
m[13'd6348]=16'h0060;
m[13'd6349]=16'h0003;
m[13'd6350]=16'h0009;
m[13'd6351]=16'ha002;
m[13'd6352]=16'h4bc1;
m[13'd6353]=16'h000a;
m[13'd6354]=16'h0009;
m[13'd6355]=16'hb009;
m[13'd6356]=16'h007b;
m[13'd6357]=16'h0301;
m[13'd6358]=16'h0009;
m[13'd6359]=16'h9b00;
m[13'd6360]=16'h0018;
m[13'd6361]=16'h4104;
m[13'd6362]=16'h0025;
m[13'd6363]=16'h4004;
m[13'd6364]=16'h004e;
m[13'd6365]=16'h0003;
m[13'd6366]=16'h0009;
m[13'd6367]=16'hb002;
m[13'd6368]=16'h4b97;
m[13'd6369]=16'h000a;
m[13'd6370]=16'h0009;
m[13'd6371]=16'hc009;
m[13'd6372]=16'h0073;
m[13'd6373]=16'h0301;
m[13'd6374]=16'h0009;
m[13'd6375]=16'h9b00;
m[13'd6376]=16'h0018;
m[13'd6377]=16'h4104;
m[13'd6378]=16'h0025;
m[13'd6379]=16'h4004;
m[13'd6380]=16'h004e;
m[13'd6381]=16'h0003;
m[13'd6382]=16'h0009;
m[13'd6383]=16'hc002;
m[13'd6384]=16'h4bae;
m[13'd6385]=16'h000a;
m[13'd6386]=16'h0009;
m[13'd6387]=16'hd009;
m[13'd6388]=16'h0073;
m[13'd6389]=16'h0301;
m[13'd6390]=16'h0009;
m[13'd6391]=16'h9b00;
m[13'd6392]=16'h0018;
m[13'd6393]=16'h4104;
m[13'd6394]=16'h0025;
m[13'd6395]=16'h4004;
m[13'd6396]=16'h004e;
m[13'd6397]=16'h0003;
m[13'd6398]=16'h0009;
m[13'd6399]=16'hd002;
m[13'd6400]=16'h4bae;
m[13'd6401]=16'h000a;
m[13'd6402]=16'h0009;
m[13'd6403]=16'he009;
m[13'd6404]=16'h0073;
m[13'd6405]=16'h0301;
m[13'd6406]=16'h0009;
m[13'd6407]=16'h9b00;
m[13'd6408]=16'h0018;
m[13'd6409]=16'h4104;
m[13'd6410]=16'h0025;
m[13'd6411]=16'h4004;
m[13'd6412]=16'h004e;
m[13'd6413]=16'h0003;
m[13'd6414]=16'h0009;
m[13'd6415]=16'he002;
m[13'd6416]=16'h4bb1;
m[13'd6417]=16'h000a;
m[13'd6418]=16'h0009;
m[13'd6419]=16'hf009;
m[13'd6420]=16'h0073;
m[13'd6421]=16'h0301;
m[13'd6422]=16'h0009;
m[13'd6423]=16'h9b00;
m[13'd6424]=16'h0018;
m[13'd6425]=16'h4104;
m[13'd6426]=16'h0025;
m[13'd6427]=16'h4004;
m[13'd6428]=16'h004e;
m[13'd6429]=16'h0003;
m[13'd6430]=16'h0009;
m[13'd6431]=16'hf002;
m[13'd6432]=16'h4bae;
m[13'd6433]=16'h010a;
m[13'd6434]=16'h0009;
m[13'd6435]=16'h0009;
m[13'd6436]=16'h0073;
m[13'd6437]=16'h0301;
m[13'd6438]=16'h0009;
m[13'd6439]=16'h9b00;
m[13'd6440]=16'h0018;
m[13'd6441]=16'h4104;
m[13'd6442]=16'h0025;
m[13'd6443]=16'h4004;
m[13'd6444]=16'h004e;
m[13'd6445]=16'h0103;
m[13'd6446]=16'h0009;
m[13'd6447]=16'h0002;
m[13'd6448]=16'h4b83;
m[13'd6449]=16'h400b;
m[13'd6450]=16'h004e;
m[13'd6451]=16'h010a;
m[13'd6452]=16'h0009;
m[13'd6453]=16'h1009;
m[13'd6454]=16'h0102;
m[13'd6455]=16'h0301;
m[13'd6456]=16'h0009;
m[13'd6457]=16'h9b00;
m[13'd6458]=16'h001b;
m[13'd6459]=16'h4002;
m[13'd6460]=16'h0010;
m[13'd6461]=16'h0003;
m[13'd6462]=16'h0016;
m[13'd6463]=16'h0905;
m[13'd6464]=16'h000a;
m[13'd6465]=16'h0906;
m[13'd6466]=16'h0007;
m[13'd6467]=16'h0004;
m[13'd6468]=16'h000a;
m[13'd6469]=16'h4104;
m[13'd6470]=16'h0095;
m[13'd6471]=16'h0003;
m[13'd6472]=16'h0009;
m[13'd6473]=16'h5002;
m[13'd6474]=16'h4a5d;
m[13'd6475]=16'h400b;
m[13'd6476]=16'h004e;
m[13'd6477]=16'h010a;
m[13'd6478]=16'h0009;
m[13'd6479]=16'h2009;
m[13'd6480]=16'h0055;
m[13'd6481]=16'h4801;
m[13'd6482]=16'h0007;
m[13'd6483]=16'h0000;
m[13'd6484]=16'h000e;
m[13'd6485]=16'h8104;
m[13'd6486]=16'h0060;
m[13'd6487]=16'h0003;
m[13'd6488]=16'h0009;
m[13'd6489]=16'h6002;
m[13'd6490]=16'h4b9d;
m[13'd6491]=16'h400b;
m[13'd6492]=16'h004e;
m[13'd6493]=16'h010a;
m[13'd6494]=16'h0009;
m[13'd6495]=16'h3009;
m[13'd6496]=16'h0073;
m[13'd6497]=16'h0301;
m[13'd6498]=16'h0009;
m[13'd6499]=16'h9b00;
m[13'd6500]=16'h0018;
m[13'd6501]=16'h4104;
m[13'd6502]=16'h0060;
m[13'd6503]=16'h0003;
m[13'd6504]=16'h0009;
m[13'd6505]=16'h7002;
m[13'd6506]=16'h4b76;
m[13'd6507]=16'h400b;
m[13'd6508]=16'h004e;
m[13'd6509]=16'h010a;
m[13'd6510]=16'h0009;
m[13'd6511]=16'h4009;
m[13'd6512]=16'h0073;
m[13'd6513]=16'h0301;
m[13'd6514]=16'h0009;
m[13'd6515]=16'h9b00;
m[13'd6516]=16'h0018;
m[13'd6517]=16'h4104;
m[13'd6518]=16'h0060;
m[13'd6519]=16'h0003;
m[13'd6520]=16'h0009;
m[13'd6521]=16'h8002;
m[13'd6522]=16'h4b73;
m[13'd6523]=16'h400b;
m[13'd6524]=16'h004e;
m[13'd6525]=16'h010a;
m[13'd6526]=16'h0009;
m[13'd6527]=16'h5009;
m[13'd6528]=16'h0073;
m[13'd6529]=16'h0301;
m[13'd6530]=16'h0009;
m[13'd6531]=16'h9b00;
m[13'd6532]=16'h0018;
m[13'd6533]=16'h4104;
m[13'd6534]=16'h0060;
m[13'd6535]=16'h0003;
m[13'd6536]=16'h0009;
m[13'd6537]=16'h9002;
m[13'd6538]=16'h4b73;
m[13'd6539]=16'h400b;
m[13'd6540]=16'h004e;
m[13'd6541]=16'h010a;
m[13'd6542]=16'h0009;
m[13'd6543]=16'h6009;
m[13'd6544]=16'h0073;
m[13'd6545]=16'h0301;
m[13'd6546]=16'h0009;
m[13'd6547]=16'h9b00;
m[13'd6548]=16'h0018;
m[13'd6549]=16'h4104;
m[13'd6550]=16'h0060;
m[13'd6551]=16'h0003;
m[13'd6552]=16'h0009;
m[13'd6553]=16'ha002;
m[13'd6554]=16'h4bc1;
m[13'd6555]=16'h010a;
m[13'd6556]=16'h0009;
m[13'd6557]=16'h7009;
m[13'd6558]=16'h007b;
m[13'd6559]=16'h0301;
m[13'd6560]=16'h0009;
m[13'd6561]=16'h9b00;
m[13'd6562]=16'h0018;
m[13'd6563]=16'h4104;
m[13'd6564]=16'h0025;
m[13'd6565]=16'h4004;
m[13'd6566]=16'h004e;
m[13'd6567]=16'h0003;
m[13'd6568]=16'h0009;
m[13'd6569]=16'hb002;
m[13'd6570]=16'h4b97;
m[13'd6571]=16'h010a;
m[13'd6572]=16'h0009;
m[13'd6573]=16'h8009;
m[13'd6574]=16'h0073;
m[13'd6575]=16'h0301;
m[13'd6576]=16'h0009;
m[13'd6577]=16'h9b00;
m[13'd6578]=16'h0018;
m[13'd6579]=16'h4104;
m[13'd6580]=16'h0025;
m[13'd6581]=16'h4004;
m[13'd6582]=16'h004e;
m[13'd6583]=16'h0003;
m[13'd6584]=16'h0009;
m[13'd6585]=16'hc002;
m[13'd6586]=16'h4bae;
m[13'd6587]=16'h010a;
m[13'd6588]=16'h0009;
m[13'd6589]=16'h9009;
m[13'd6590]=16'h0073;
m[13'd6591]=16'h0301;
m[13'd6592]=16'h0009;
m[13'd6593]=16'h9b00;
m[13'd6594]=16'h0018;
m[13'd6595]=16'h4104;
m[13'd6596]=16'h0025;
m[13'd6597]=16'h4004;
m[13'd6598]=16'h004e;
m[13'd6599]=16'h0003;
m[13'd6600]=16'h0009;
m[13'd6601]=16'hd002;
m[13'd6602]=16'h4bae;
m[13'd6603]=16'h010a;
m[13'd6604]=16'h0009;
m[13'd6605]=16'ha009;
m[13'd6606]=16'h0073;
m[13'd6607]=16'h0301;
m[13'd6608]=16'h0009;
m[13'd6609]=16'h9b00;
m[13'd6610]=16'h0018;
m[13'd6611]=16'h4104;
m[13'd6612]=16'h0025;
m[13'd6613]=16'h4004;
m[13'd6614]=16'h004e;
m[13'd6615]=16'h0003;
m[13'd6616]=16'h0009;
m[13'd6617]=16'he002;
m[13'd6618]=16'h4bb1;
m[13'd6619]=16'h010a;
m[13'd6620]=16'h0009;
m[13'd6621]=16'hb009;
m[13'd6622]=16'h0073;
m[13'd6623]=16'h0301;
m[13'd6624]=16'h0009;
m[13'd6625]=16'h9b00;
m[13'd6626]=16'h0018;
m[13'd6627]=16'h4104;
m[13'd6628]=16'h0025;
m[13'd6629]=16'h4004;
m[13'd6630]=16'h004e;
m[13'd6631]=16'h0003;
m[13'd6632]=16'h0009;
m[13'd6633]=16'hf002;
m[13'd6634]=16'h4bae;
m[13'd6635]=16'h010a;
m[13'd6636]=16'h0009;
m[13'd6637]=16'hc009;
m[13'd6638]=16'h0073;
m[13'd6639]=16'h0301;
m[13'd6640]=16'h0009;
m[13'd6641]=16'h9b00;
m[13'd6642]=16'h0018;
m[13'd6643]=16'h4104;
m[13'd6644]=16'h0025;
m[13'd6645]=16'h4004;
m[13'd6646]=16'h004e;
m[13'd6647]=16'h0103;
m[13'd6648]=16'h0009;
m[13'd6649]=16'h0002;
m[13'd6650]=16'h4c0b;
m[13'd6651]=16'h0108;
m[13'd6652]=16'h0009;
m[13'd6653]=16'h2307;
m[13'd6654]=16'h001b;
m[13'd6655]=16'h4009;
m[13'd6656]=16'h0010;
m[13'd6657]=16'h000a;
m[13'd6658]=16'h0016;
m[13'd6659]=16'h090c;
m[13'd6660]=16'h000a;
m[13'd6661]=16'h090d;
m[13'd6662]=16'h0007;
m[13'd6663]=16'h000b;
m[13'd6664]=16'h000a;
m[13'd6665]=16'h410b;
m[13'd6666]=16'h0095;
m[13'd6667]=16'h000a;
m[13'd6668]=16'h0009;
m[13'd6669]=16'h5009;
m[13'd6670]=16'h010f;
m[13'd6671]=16'h0301;
m[13'd6672]=16'h0009;
m[13'd6673]=16'h9b00;
m[13'd6674]=16'h001b;
m[13'd6675]=16'h4002;
m[13'd6676]=16'h0010;
m[13'd6677]=16'h0003;
m[13'd6678]=16'h0016;
m[13'd6679]=16'h0905;
m[13'd6680]=16'h000a;
m[13'd6681]=16'h0906;
m[13'd6682]=16'h0007;
m[13'd6683]=16'h0004;
m[13'd6684]=16'h000a;
m[13'd6685]=16'h4104;
m[13'd6686]=16'h008d;
m[13'd6687]=16'h0003;
m[13'd6688]=16'h0009;
m[13'd6689]=16'h5002;
m[13'd6690]=16'h4927;
m[13'd6691]=16'h810b;
m[13'd6692]=16'h002b;
m[13'd6693]=16'h3108;
m[13'd6694]=16'h0007;
m[13'd6695]=16'h0007;
m[13'd6696]=16'h0060;
m[13'd6697]=16'h000a;
m[13'd6698]=16'h0009;
m[13'd6699]=16'h6009;
m[13'd6700]=16'h0055;
m[13'd6701]=16'h4801;
m[13'd6702]=16'h0007;
m[13'd6703]=16'h0000;
m[13'd6704]=16'h000e;
m[13'd6705]=16'h8104;
m[13'd6706]=16'h0058;
m[13'd6707]=16'h0003;
m[13'd6708]=16'h0009;
m[13'd6709]=16'h6002;
m[13'd6710]=16'h4b60;
m[13'd6711]=16'h110b;
m[13'd6712]=16'h002b;
m[13'd6713]=16'h1108;
m[13'd6714]=16'h0007;
m[13'd6715]=16'h0007;
m[13'd6716]=16'h0060;
m[13'd6717]=16'h000a;
m[13'd6718]=16'h0009;
m[13'd6719]=16'h7009;
m[13'd6720]=16'h0073;
m[13'd6721]=16'h0301;
m[13'd6722]=16'h0009;
m[13'd6723]=16'h9b00;
m[13'd6724]=16'h0018;
m[13'd6725]=16'h4104;
m[13'd6726]=16'h0058;
m[13'd6727]=16'h0003;
m[13'd6728]=16'h0009;
m[13'd6729]=16'h7002;
m[13'd6730]=16'h4b39;
m[13'd6731]=16'h800b;
m[13'd6732]=16'h002b;
m[13'd6733]=16'h0808;
m[13'd6734]=16'h0007;
m[13'd6735]=16'h0007;
m[13'd6736]=16'h0060;
m[13'd6737]=16'h000a;
m[13'd6738]=16'h0009;
m[13'd6739]=16'h8009;
m[13'd6740]=16'h0073;
m[13'd6741]=16'h0301;
m[13'd6742]=16'h0009;
m[13'd6743]=16'h9b00;
m[13'd6744]=16'h0018;
m[13'd6745]=16'h4104;
m[13'd6746]=16'h0058;
m[13'd6747]=16'h0003;
m[13'd6748]=16'h0009;
m[13'd6749]=16'h8002;
m[13'd6750]=16'h4b39;
m[13'd6751]=16'h400b;
m[13'd6752]=16'h002b;
m[13'd6753]=16'h1608;
m[13'd6754]=16'h0007;
m[13'd6755]=16'h0007;
m[13'd6756]=16'h0060;
m[13'd6757]=16'h000a;
m[13'd6758]=16'h0009;
m[13'd6759]=16'h9009;
m[13'd6760]=16'h0073;
m[13'd6761]=16'h0301;
m[13'd6762]=16'h0009;
m[13'd6763]=16'h9b00;
m[13'd6764]=16'h0018;
m[13'd6765]=16'h4104;
m[13'd6766]=16'h0058;
m[13'd6767]=16'h0003;
m[13'd6768]=16'h0009;
m[13'd6769]=16'h9002;
m[13'd6770]=16'h4b36;
m[13'd6771]=16'h800b;
m[13'd6772]=16'h002b;
m[13'd6773]=16'h0508;
m[13'd6774]=16'h0007;
m[13'd6775]=16'h0007;
m[13'd6776]=16'h0060;
m[13'd6777]=16'h000a;
m[13'd6778]=16'h0009;
m[13'd6779]=16'ha009;
m[13'd6780]=16'h0073;
m[13'd6781]=16'h0301;
m[13'd6782]=16'h0009;
m[13'd6783]=16'h9b00;
m[13'd6784]=16'h0018;
m[13'd6785]=16'h4104;
m[13'd6786]=16'h0058;
m[13'd6787]=16'h0003;
m[13'd6788]=16'h0009;
m[13'd6789]=16'ha002;
m[13'd6790]=16'h4b49;
m[13'd6791]=16'h800b;
m[13'd6792]=16'h002b;
m[13'd6793]=16'h0408;
m[13'd6794]=16'h0007;
m[13'd6795]=16'h0007;
m[13'd6796]=16'h0025;
m[13'd6797]=16'h400b;
m[13'd6798]=16'h004e;
m[13'd6799]=16'h000a;
m[13'd6800]=16'h0009;
m[13'd6801]=16'hb009;
m[13'd6802]=16'h0102;
m[13'd6803]=16'h0401;
m[13'd6804]=16'h0009;
m[13'd6805]=16'h4900;
m[13'd6806]=16'h001b;
m[13'd6807]=16'h4002;
m[13'd6808]=16'h0010;
m[13'd6809]=16'h0003;
m[13'd6810]=16'h0016;
m[13'd6811]=16'h0905;
m[13'd6812]=16'h000a;
m[13'd6813]=16'h0906;
m[13'd6814]=16'h0007;
m[13'd6815]=16'h0004;
m[13'd6816]=16'h000a;
m[13'd6817]=16'h4104;
m[13'd6818]=16'h008d;
m[13'd6819]=16'h0003;
m[13'd6820]=16'h0009;
m[13'd6821]=16'h5002;
m[13'd6822]=16'h4a0e;
m[13'd6823]=16'h800b;
m[13'd6824]=16'h002b;
m[13'd6825]=16'h0308;
m[13'd6826]=16'h0007;
m[13'd6827]=16'h0007;
m[13'd6828]=16'h0025;
m[13'd6829]=16'h400b;
m[13'd6830]=16'h004e;
m[13'd6831]=16'h000a;
m[13'd6832]=16'h0009;
m[13'd6833]=16'hc009;
m[13'd6834]=16'h0055;
m[13'd6835]=16'h4801;
m[13'd6836]=16'h0007;
m[13'd6837]=16'h0000;
m[13'd6838]=16'h000e;
m[13'd6839]=16'h8104;
m[13'd6840]=16'h0058;
m[13'd6841]=16'h0003;
m[13'd6842]=16'h0009;
m[13'd6843]=16'h6002;
m[13'd6844]=16'h4b4e;
m[13'd6845]=16'h800b;
m[13'd6846]=16'h002b;
m[13'd6847]=16'h0308;
m[13'd6848]=16'h0007;
m[13'd6849]=16'h0007;
m[13'd6850]=16'h0025;
m[13'd6851]=16'h400b;
m[13'd6852]=16'h004e;
m[13'd6853]=16'h000a;
m[13'd6854]=16'h0009;
m[13'd6855]=16'hd009;
m[13'd6856]=16'h0073;
m[13'd6857]=16'h0401;
m[13'd6858]=16'h0009;
m[13'd6859]=16'h4900;
m[13'd6860]=16'h0018;
m[13'd6861]=16'h4104;
m[13'd6862]=16'h0058;
m[13'd6863]=16'h0003;
m[13'd6864]=16'h0009;
m[13'd6865]=16'h7002;
m[13'd6866]=16'h4b24;
m[13'd6867]=16'h100b;
m[13'd6868]=16'h002b;
m[13'd6869]=16'h1208;
m[13'd6870]=16'h0007;
m[13'd6871]=16'h0007;
m[13'd6872]=16'h0025;
m[13'd6873]=16'h400b;
m[13'd6874]=16'h004e;
m[13'd6875]=16'h000a;
m[13'd6876]=16'h0009;
m[13'd6877]=16'he009;
m[13'd6878]=16'h0073;
m[13'd6879]=16'h0401;
m[13'd6880]=16'h0009;
m[13'd6881]=16'h4900;
m[13'd6882]=16'h0018;
m[13'd6883]=16'h4104;
m[13'd6884]=16'h0058;
m[13'd6885]=16'h0003;
m[13'd6886]=16'h0009;
m[13'd6887]=16'h8002;
m[13'd6888]=16'h4b27;
m[13'd6889]=16'h100b;
m[13'd6890]=16'h002b;
m[13'd6891]=16'h1208;
m[13'd6892]=16'h0007;
m[13'd6893]=16'h0007;
m[13'd6894]=16'h0025;
m[13'd6895]=16'h400b;
m[13'd6896]=16'h004e;
m[13'd6897]=16'h000a;
m[13'd6898]=16'h0009;
m[13'd6899]=16'hf009;
m[13'd6900]=16'h0073;
m[13'd6901]=16'h0401;
m[13'd6902]=16'h0009;
m[13'd6903]=16'h4900;
m[13'd6904]=16'h0018;
m[13'd6905]=16'h4104;
m[13'd6906]=16'h0058;
m[13'd6907]=16'h0003;
m[13'd6908]=16'h0009;
m[13'd6909]=16'h9002;
m[13'd6910]=16'h4b24;
m[13'd6911]=16'h100b;
m[13'd6912]=16'h002b;
m[13'd6913]=16'h1108;
m[13'd6914]=16'h0007;
m[13'd6915]=16'h0007;
m[13'd6916]=16'h0025;
m[13'd6917]=16'h400b;
m[13'd6918]=16'h004e;
m[13'd6919]=16'h010a;
m[13'd6920]=16'h0009;
m[13'd6921]=16'h0009;
m[13'd6922]=16'h0073;
m[13'd6923]=16'h0401;
m[13'd6924]=16'h0009;
m[13'd6925]=16'h4900;
m[13'd6926]=16'h0018;
m[13'd6927]=16'h4104;
m[13'd6928]=16'h0058;
m[13'd6929]=16'h0003;
m[13'd6930]=16'h0009;
m[13'd6931]=16'ha002;
m[13'd6932]=16'h4bae;
m[13'd6933]=16'h0808;
m[13'd6934]=16'h0009;
m[13'd6935]=16'h9307;
m[13'd6936]=16'h001b;
m[13'd6937]=16'h4009;
m[13'd6938]=16'h0010;
m[13'd6939]=16'h000a;
m[13'd6940]=16'h0016;
m[13'd6941]=16'h090c;
m[13'd6942]=16'h000a;
m[13'd6943]=16'h090d;
m[13'd6944]=16'h0007;
m[13'd6945]=16'h000b;
m[13'd6946]=16'h000a;
m[13'd6947]=16'h410b;
m[13'd6948]=16'h0095;
m[13'd6949]=16'h000a;
m[13'd6950]=16'h0009;
m[13'd6951]=16'h5009;
m[13'd6952]=16'h010f;
m[13'd6953]=16'h0301;
m[13'd6954]=16'h0009;
m[13'd6955]=16'h9b00;
m[13'd6956]=16'h001b;
m[13'd6957]=16'h4002;
m[13'd6958]=16'h0010;
m[13'd6959]=16'h0003;
m[13'd6960]=16'h0016;
m[13'd6961]=16'h0905;
m[13'd6962]=16'h000a;
m[13'd6963]=16'h0906;
m[13'd6964]=16'h0007;
m[13'd6965]=16'h0004;
m[13'd6966]=16'h000a;
m[13'd6967]=16'h4104;
m[13'd6968]=16'h0095;
m[13'd6969]=16'h0003;
m[13'd6970]=16'h0009;
m[13'd6971]=16'h5002;
m[13'd6972]=16'h4963;
m[13'd6973]=16'h000a;
m[13'd6974]=16'h0009;
m[13'd6975]=16'h6009;
m[13'd6976]=16'h0055;
m[13'd6977]=16'h4801;
m[13'd6978]=16'h0007;
m[13'd6979]=16'h0000;
m[13'd6980]=16'h000e;
m[13'd6981]=16'h8104;
m[13'd6982]=16'h0060;
m[13'd6983]=16'h0003;
m[13'd6984]=16'h0009;
m[13'd6985]=16'h6002;
m[13'd6986]=16'h4bed;
m[13'd6987]=16'h000a;
m[13'd6988]=16'h0009;
m[13'd6989]=16'h7009;
m[13'd6990]=16'h0073;
m[13'd6991]=16'h0301;
m[13'd6992]=16'h0009;
m[13'd6993]=16'h9b00;
m[13'd6994]=16'h0018;
m[13'd6995]=16'h4104;
m[13'd6996]=16'h0060;
m[13'd6997]=16'h0003;
m[13'd6998]=16'h0009;
m[13'd6999]=16'h7002;
m[13'd7000]=16'h4bc0;
m[13'd7001]=16'h000a;
m[13'd7002]=16'h0009;
m[13'd7003]=16'h8009;
m[13'd7004]=16'h0073;
m[13'd7005]=16'h0301;
m[13'd7006]=16'h0009;
m[13'd7007]=16'h9b00;
m[13'd7008]=16'h0018;
m[13'd7009]=16'h4104;
m[13'd7010]=16'h0060;
m[13'd7011]=16'h0003;
m[13'd7012]=16'h0009;
m[13'd7013]=16'h8002;
m[13'd7014]=16'h4bc3;
m[13'd7015]=16'h000a;
m[13'd7016]=16'h0009;
m[13'd7017]=16'h9009;
m[13'd7018]=16'h0073;
m[13'd7019]=16'h0301;
m[13'd7020]=16'h0009;
m[13'd7021]=16'h9b00;
m[13'd7022]=16'h0018;
m[13'd7023]=16'h4104;
m[13'd7024]=16'h0060;
m[13'd7025]=16'h0003;
m[13'd7026]=16'h0009;
m[13'd7027]=16'h9002;
m[13'd7028]=16'h4bc3;
m[13'd7029]=16'h000a;
m[13'd7030]=16'h0009;
m[13'd7031]=16'ha009;
m[13'd7032]=16'h0073;
m[13'd7033]=16'h0301;
m[13'd7034]=16'h0009;
m[13'd7035]=16'h9b00;
m[13'd7036]=16'h0018;
m[13'd7037]=16'h4104;
m[13'd7038]=16'h0060;
m[13'd7039]=16'h0003;
m[13'd7040]=16'h0009;
m[13'd7041]=16'ha002;
m[13'd7042]=16'h4b95;
m[13'd7043]=16'h400b;
m[13'd7044]=16'h004e;
m[13'd7045]=16'h000a;
m[13'd7046]=16'h0009;
m[13'd7047]=16'hb009;
m[13'd7048]=16'h007b;
m[13'd7049]=16'h0301;
m[13'd7050]=16'h0009;
m[13'd7051]=16'h9b00;
m[13'd7052]=16'h0018;
m[13'd7053]=16'h4104;
m[13'd7054]=16'h0025;
m[13'd7055]=16'h4004;
m[13'd7056]=16'h004e;
m[13'd7057]=16'h0003;
m[13'd7058]=16'h0009;
m[13'd7059]=16'hb002;
m[13'd7060]=16'h4b4a;
m[13'd7061]=16'h400b;
m[13'd7062]=16'h004e;
m[13'd7063]=16'h000a;
m[13'd7064]=16'h0009;
m[13'd7065]=16'hc009;
m[13'd7066]=16'h0073;
m[13'd7067]=16'h0301;
m[13'd7068]=16'h0009;
m[13'd7069]=16'h9b00;
m[13'd7070]=16'h0018;
m[13'd7071]=16'h4104;
m[13'd7072]=16'h0025;
m[13'd7073]=16'h4004;
m[13'd7074]=16'h004e;
m[13'd7075]=16'h0003;
m[13'd7076]=16'h0009;
m[13'd7077]=16'hc002;
m[13'd7078]=16'h4b61;
m[13'd7079]=16'h400b;
m[13'd7080]=16'h004e;
m[13'd7081]=16'h000a;
m[13'd7082]=16'h0009;
m[13'd7083]=16'hd009;
m[13'd7084]=16'h0073;
m[13'd7085]=16'h0301;
m[13'd7086]=16'h0009;
m[13'd7087]=16'h9b00;
m[13'd7088]=16'h0018;
m[13'd7089]=16'h4104;
m[13'd7090]=16'h0025;
m[13'd7091]=16'h4004;
m[13'd7092]=16'h004e;
m[13'd7093]=16'h0003;
m[13'd7094]=16'h0009;
m[13'd7095]=16'hd002;
m[13'd7096]=16'h4b61;
m[13'd7097]=16'h400b;
m[13'd7098]=16'h004e;
m[13'd7099]=16'h000a;
m[13'd7100]=16'h0009;
m[13'd7101]=16'he009;
m[13'd7102]=16'h0073;
m[13'd7103]=16'h0301;
m[13'd7104]=16'h0009;
m[13'd7105]=16'h9b00;
m[13'd7106]=16'h0018;
m[13'd7107]=16'h4104;
m[13'd7108]=16'h0025;
m[13'd7109]=16'h4004;
m[13'd7110]=16'h004e;
m[13'd7111]=16'h0003;
m[13'd7112]=16'h0009;
m[13'd7113]=16'he002;
m[13'd7114]=16'h4b61;
m[13'd7115]=16'h400b;
m[13'd7116]=16'h004e;
m[13'd7117]=16'h000a;
m[13'd7118]=16'h0009;
m[13'd7119]=16'hf009;
m[13'd7120]=16'h0073;
m[13'd7121]=16'h0301;
m[13'd7122]=16'h0009;
m[13'd7123]=16'h9b00;
m[13'd7124]=16'h0018;
m[13'd7125]=16'h4104;
m[13'd7126]=16'h0025;
m[13'd7127]=16'h4004;
m[13'd7128]=16'h004e;
m[13'd7129]=16'h0003;
m[13'd7130]=16'h0009;
m[13'd7131]=16'hf002;
m[13'd7132]=16'h4b61;
m[13'd7133]=16'h400b;
m[13'd7134]=16'h004e;
m[13'd7135]=16'h010a;
m[13'd7136]=16'h0009;
m[13'd7137]=16'h0009;
m[13'd7138]=16'h0073;
m[13'd7139]=16'h0301;
m[13'd7140]=16'h0009;
m[13'd7141]=16'h9b00;
m[13'd7142]=16'h0018;
m[13'd7143]=16'h4104;
m[13'd7144]=16'h0025;
m[13'd7145]=16'h4004;
m[13'd7146]=16'h004e;
m[13'd7147]=16'h0103;
m[13'd7148]=16'h0009;
m[13'd7149]=16'h0002;
m[13'd7150]=16'h4be3;
m[13'd7151]=16'h0908;
m[13'd7152]=16'h0009;
m[13'd7153]=16'h9f07;
m[13'd7154]=16'h001b;
m[13'd7155]=16'h4009;
m[13'd7156]=16'h0010;
m[13'd7157]=16'h000a;
m[13'd7158]=16'h0016;
m[13'd7159]=16'h090c;
m[13'd7160]=16'h000a;
m[13'd7161]=16'h090d;
m[13'd7162]=16'h0007;
m[13'd7163]=16'h000b;
m[13'd7164]=16'h000a;
m[13'd7165]=16'h410b;
m[13'd7166]=16'h0095;
m[13'd7167]=16'h000a;
m[13'd7168]=16'h0009;
m[13'd7169]=16'h5009;
m[13'd7170]=16'h010f;
m[13'd7171]=16'h0401;
m[13'd7172]=16'h0009;
m[13'd7173]=16'hd000;
m[13'd7174]=16'h001b;
m[13'd7175]=16'h4002;
m[13'd7176]=16'h0010;
m[13'd7177]=16'h0003;
m[13'd7178]=16'h0016;
m[13'd7179]=16'h0905;
m[13'd7180]=16'h000a;
m[13'd7181]=16'h0906;
m[13'd7182]=16'h0007;
m[13'd7183]=16'h0004;
m[13'd7184]=16'h000a;
m[13'd7185]=16'h4104;
m[13'd7186]=16'h008d;
m[13'd7187]=16'h0003;
m[13'd7188]=16'h0009;
m[13'd7189]=16'h5002;
m[13'd7190]=16'h4975;
m[13'd7191]=16'h000a;
m[13'd7192]=16'h0009;
m[13'd7193]=16'h6009;
m[13'd7194]=16'h0055;
m[13'd7195]=16'h4801;
m[13'd7196]=16'h0007;
m[13'd7197]=16'h0000;
m[13'd7198]=16'h000e;
m[13'd7199]=16'h8104;
m[13'd7200]=16'h0058;
m[13'd7201]=16'h0003;
m[13'd7202]=16'h0009;
m[13'd7203]=16'h6002;
m[13'd7204]=16'h4bf3;
m[13'd7205]=16'h000a;
m[13'd7206]=16'h0009;
m[13'd7207]=16'h7009;
m[13'd7208]=16'h0073;
m[13'd7209]=16'h0401;
m[13'd7210]=16'h0009;
m[13'd7211]=16'hd000;
m[13'd7212]=16'h0018;
m[13'd7213]=16'h4104;
m[13'd7214]=16'h0058;
m[13'd7215]=16'h0003;
m[13'd7216]=16'h0009;
m[13'd7217]=16'h7002;
m[13'd7218]=16'h4bc9;
m[13'd7219]=16'h000a;
m[13'd7220]=16'h0009;
m[13'd7221]=16'h8009;
m[13'd7222]=16'h0073;
m[13'd7223]=16'h0401;
m[13'd7224]=16'h0009;
m[13'd7225]=16'hd000;
m[13'd7226]=16'h0018;
m[13'd7227]=16'h4104;
m[13'd7228]=16'h0058;
m[13'd7229]=16'h0003;
m[13'd7230]=16'h0009;
m[13'd7231]=16'h8002;
m[13'd7232]=16'h4bcc;
m[13'd7233]=16'h000a;
m[13'd7234]=16'h0009;
m[13'd7235]=16'h9009;
m[13'd7236]=16'h0073;
m[13'd7237]=16'h0401;
m[13'd7238]=16'h0009;
m[13'd7239]=16'hd000;
m[13'd7240]=16'h0018;
m[13'd7241]=16'h4104;
m[13'd7242]=16'h0058;
m[13'd7243]=16'h0003;
m[13'd7244]=16'h0009;
m[13'd7245]=16'h9002;
m[13'd7246]=16'h4bc9;
m[13'd7247]=16'h000a;
m[13'd7248]=16'h0009;
m[13'd7249]=16'ha009;
m[13'd7250]=16'h0073;
m[13'd7251]=16'h0401;
m[13'd7252]=16'h0009;
m[13'd7253]=16'hd000;
m[13'd7254]=16'h0018;
m[13'd7255]=16'h4104;
m[13'd7256]=16'h0058;
m[13'd7257]=16'h0003;
m[13'd7258]=16'h0009;
m[13'd7259]=16'ha002;
m[13'd7260]=16'h4b9e;
m[13'd7261]=16'h400b;
m[13'd7262]=16'h004e;
m[13'd7263]=16'h000a;
m[13'd7264]=16'h0009;
m[13'd7265]=16'hb009;
m[13'd7266]=16'h0102;
m[13'd7267]=16'h0501;
m[13'd7268]=16'h0009;
m[13'd7269]=16'h1900;
m[13'd7270]=16'h001b;
m[13'd7271]=16'h4002;
m[13'd7272]=16'h0010;
m[13'd7273]=16'h0003;
m[13'd7274]=16'h0016;
m[13'd7275]=16'h0905;
m[13'd7276]=16'h000a;
m[13'd7277]=16'h0906;
m[13'd7278]=16'h0007;
m[13'd7279]=16'h0004;
m[13'd7280]=16'h000a;
m[13'd7281]=16'h4104;
m[13'd7282]=16'h008d;
m[13'd7283]=16'h0003;
m[13'd7284]=16'h0009;
m[13'd7285]=16'h5002;
m[13'd7286]=16'h4a66;
m[13'd7287]=16'h400b;
m[13'd7288]=16'h004e;
m[13'd7289]=16'h000a;
m[13'd7290]=16'h0009;
m[13'd7291]=16'hc009;
m[13'd7292]=16'h0055;
m[13'd7293]=16'h4801;
m[13'd7294]=16'h0007;
m[13'd7295]=16'h0000;
m[13'd7296]=16'h000e;
m[13'd7297]=16'h8104;
m[13'd7298]=16'h0058;
m[13'd7299]=16'h0003;
m[13'd7300]=16'h0009;
m[13'd7301]=16'h6002;
m[13'd7302]=16'h4ba6;
m[13'd7303]=16'h400b;
m[13'd7304]=16'h004e;
m[13'd7305]=16'h000a;
m[13'd7306]=16'h0009;
m[13'd7307]=16'hd009;
m[13'd7308]=16'h0073;
m[13'd7309]=16'h0501;
m[13'd7310]=16'h0009;
m[13'd7311]=16'h1900;
m[13'd7312]=16'h0018;
m[13'd7313]=16'h4104;
m[13'd7314]=16'h0058;
m[13'd7315]=16'h0003;
m[13'd7316]=16'h0009;
m[13'd7317]=16'h7002;
m[13'd7318]=16'h4b7c;
m[13'd7319]=16'h400b;
m[13'd7320]=16'h004e;
m[13'd7321]=16'h000a;
m[13'd7322]=16'h0009;
m[13'd7323]=16'he009;
m[13'd7324]=16'h0073;
m[13'd7325]=16'h0501;
m[13'd7326]=16'h0009;
m[13'd7327]=16'h1900;
m[13'd7328]=16'h0018;
m[13'd7329]=16'h4104;
m[13'd7330]=16'h0058;
m[13'd7331]=16'h0003;
m[13'd7332]=16'h0009;
m[13'd7333]=16'h8002;
m[13'd7334]=16'h4b7c;
m[13'd7335]=16'h400b;
m[13'd7336]=16'h004e;
m[13'd7337]=16'h000a;
m[13'd7338]=16'h0009;
m[13'd7339]=16'hf009;
m[13'd7340]=16'h0073;
m[13'd7341]=16'h0501;
m[13'd7342]=16'h0009;
m[13'd7343]=16'h1900;
m[13'd7344]=16'h0018;
m[13'd7345]=16'h4104;
m[13'd7346]=16'h0058;
m[13'd7347]=16'h0003;
m[13'd7348]=16'h0009;
m[13'd7349]=16'h9002;
m[13'd7350]=16'h4b7c;
m[13'd7351]=16'h400b;
m[13'd7352]=16'h004e;
m[13'd7353]=16'h010a;
m[13'd7354]=16'h0009;
m[13'd7355]=16'h0009;
m[13'd7356]=16'h0073;
m[13'd7357]=16'h0501;
m[13'd7358]=16'h0009;
m[13'd7359]=16'h1900;
m[13'd7360]=16'h0018;
m[13'd7361]=16'h4104;
m[13'd7362]=16'h0058;
m[13'd7363]=16'h0003;
m[13'd7364]=16'h0009;
m[13'd7365]=16'ha002;
m[13'd7366]=16'h4bc7;
m[13'd7367]=16'h010a;
m[13'd7368]=16'h0009;
m[13'd7369]=16'h1009;
m[13'd7370]=16'h0102;
m[13'd7371]=16'h0501;
m[13'd7372]=16'h0009;
m[13'd7373]=16'h6700;
m[13'd7374]=16'h001b;
m[13'd7375]=16'h4002;
m[13'd7376]=16'h0010;
m[13'd7377]=16'h0003;
m[13'd7378]=16'h0016;
m[13'd7379]=16'h0905;
m[13'd7380]=16'h000a;
m[13'd7381]=16'h0906;
m[13'd7382]=16'h0007;
m[13'd7383]=16'h0004;
m[13'd7384]=16'h000a;
m[13'd7385]=16'h4104;
m[13'd7386]=16'h008d;
m[13'd7387]=16'h0003;
m[13'd7388]=16'h0009;
m[13'd7389]=16'h5002;
m[13'd7390]=16'h4ab0;
m[13'd7391]=16'h010a;
m[13'd7392]=16'h0009;
m[13'd7393]=16'h2009;
m[13'd7394]=16'h0055;
m[13'd7395]=16'h4801;
m[13'd7396]=16'h0007;
m[13'd7397]=16'h0000;
m[13'd7398]=16'h000e;
m[13'd7399]=16'h8104;
m[13'd7400]=16'h0058;
m[13'd7401]=16'h0003;
m[13'd7402]=16'h0009;
m[13'd7403]=16'h6002;
m[13'd7404]=16'h4bf6;
m[13'd7405]=16'h010a;
m[13'd7406]=16'h0009;
m[13'd7407]=16'h3009;
m[13'd7408]=16'h0073;
m[13'd7409]=16'h0501;
m[13'd7410]=16'h0009;
m[13'd7411]=16'h6700;
m[13'd7412]=16'h0018;
m[13'd7413]=16'h4104;
m[13'd7414]=16'h0058;
m[13'd7415]=16'h0003;
m[13'd7416]=16'h0009;
m[13'd7417]=16'h7002;
m[13'd7418]=16'h4bc9;
m[13'd7419]=16'h010a;
m[13'd7420]=16'h0009;
m[13'd7421]=16'h4009;
m[13'd7422]=16'h0073;
m[13'd7423]=16'h0501;
m[13'd7424]=16'h0009;
m[13'd7425]=16'h6700;
m[13'd7426]=16'h0018;
m[13'd7427]=16'h4104;
m[13'd7428]=16'h0058;
m[13'd7429]=16'h0003;
m[13'd7430]=16'h0009;
m[13'd7431]=16'h8002;
m[13'd7432]=16'h4bc9;
m[13'd7433]=16'h010a;
m[13'd7434]=16'h0009;
m[13'd7435]=16'h5009;
m[13'd7436]=16'h0073;
m[13'd7437]=16'h0501;
m[13'd7438]=16'h0009;
m[13'd7439]=16'h6700;
m[13'd7440]=16'h0018;
m[13'd7441]=16'h4104;
m[13'd7442]=16'h0058;
m[13'd7443]=16'h0003;
m[13'd7444]=16'h0009;
m[13'd7445]=16'h9002;
m[13'd7446]=16'h4bcc;
m[13'd7447]=16'h010a;
m[13'd7448]=16'h0009;
m[13'd7449]=16'h6009;
m[13'd7450]=16'h0073;
m[13'd7451]=16'h0501;
m[13'd7452]=16'h0009;
m[13'd7453]=16'h6700;
m[13'd7454]=16'h0018;
m[13'd7455]=16'h4104;
m[13'd7456]=16'h0058;
m[13'd7457]=16'h0003;
m[13'd7458]=16'h0009;
m[13'd7459]=16'ha002;
m[13'd7460]=16'h4c10;
m[13'd7461]=16'h0808;
m[13'd7462]=16'h0009;
m[13'd7463]=16'h9307;
m[13'd7464]=16'h001b;
m[13'd7465]=16'h4009;
m[13'd7466]=16'h0010;
m[13'd7467]=16'h000a;
m[13'd7468]=16'h0016;
m[13'd7469]=16'h090c;
m[13'd7470]=16'h000a;
m[13'd7471]=16'h090d;
m[13'd7472]=16'h0007;
m[13'd7473]=16'h000b;
m[13'd7474]=16'h000a;
m[13'd7475]=16'h410b;
m[13'd7476]=16'h008d;
m[13'd7477]=16'h000a;
m[13'd7478]=16'h0009;
m[13'd7479]=16'h5009;
m[13'd7480]=16'h0110;
m[13'd7481]=16'h0601;
m[13'd7482]=16'h0009;
m[13'd7483]=16'h6c00;
m[13'd7484]=16'h001b;
m[13'd7485]=16'h4002;
m[13'd7486]=16'h0010;
m[13'd7487]=16'h0003;
m[13'd7488]=16'h0016;
m[13'd7489]=16'h0905;
m[13'd7490]=16'h000a;
m[13'd7491]=16'h0906;
m[13'd7492]=16'h0007;
m[13'd7493]=16'h0004;
m[13'd7494]=16'h000a;
m[13'd7495]=16'h4104;
m[13'd7496]=16'h0095;
m[13'd7497]=16'h0003;
m[13'd7498]=16'h0009;
m[13'd7499]=16'h5002;
m[13'd7500]=16'h496a;
m[13'd7501]=16'h000a;
m[13'd7502]=16'h0009;
m[13'd7503]=16'h6009;
m[13'd7504]=16'h0055;
m[13'd7505]=16'h4801;
m[13'd7506]=16'h0007;
m[13'd7507]=16'h0000;
m[13'd7508]=16'h000e;
m[13'd7509]=16'h8104;
m[13'd7510]=16'h0060;
m[13'd7511]=16'h0003;
m[13'd7512]=16'h0009;
m[13'd7513]=16'h6002;
m[13'd7514]=16'h4bee;
m[13'd7515]=16'h000a;
m[13'd7516]=16'h0009;
m[13'd7517]=16'h7009;
m[13'd7518]=16'h0074;
m[13'd7519]=16'h0601;
m[13'd7520]=16'h0009;
m[13'd7521]=16'h6c00;
m[13'd7522]=16'h0018;
m[13'd7523]=16'h4104;
m[13'd7524]=16'h0060;
m[13'd7525]=16'h0003;
m[13'd7526]=16'h0009;
m[13'd7527]=16'h7002;
m[13'd7528]=16'h4bc1;
m[13'd7529]=16'h000a;
m[13'd7530]=16'h0009;
m[13'd7531]=16'h8009;
m[13'd7532]=16'h0074;
m[13'd7533]=16'h0601;
m[13'd7534]=16'h0009;
m[13'd7535]=16'h6c00;
m[13'd7536]=16'h0018;
m[13'd7537]=16'h4104;
m[13'd7538]=16'h0060;
m[13'd7539]=16'h0003;
m[13'd7540]=16'h0009;
m[13'd7541]=16'h8002;
m[13'd7542]=16'h4bc1;
m[13'd7543]=16'h000a;
m[13'd7544]=16'h0009;
m[13'd7545]=16'h9009;
m[13'd7546]=16'h0074;
m[13'd7547]=16'h0601;
m[13'd7548]=16'h0009;
m[13'd7549]=16'h6c00;
m[13'd7550]=16'h0018;
m[13'd7551]=16'h4104;
m[13'd7552]=16'h0060;
m[13'd7553]=16'h0003;
m[13'd7554]=16'h0009;
m[13'd7555]=16'h9002;
m[13'd7556]=16'h4bc1;
m[13'd7557]=16'h000a;
m[13'd7558]=16'h0009;
m[13'd7559]=16'ha009;
m[13'd7560]=16'h0074;
m[13'd7561]=16'h0601;
m[13'd7562]=16'h0009;
m[13'd7563]=16'h6c00;
m[13'd7564]=16'h0018;
m[13'd7565]=16'h4104;
m[13'd7566]=16'h0060;
m[13'd7567]=16'h0003;
m[13'd7568]=16'h0009;
m[13'd7569]=16'ha002;
m[13'd7570]=16'h4c26;
m[13'd7571]=16'h0108;
m[13'd7572]=16'h0009;
m[13'd7573]=16'h2307;
m[13'd7574]=16'h001b;
m[13'd7575]=16'h4009;
m[13'd7576]=16'h0010;
m[13'd7577]=16'h000a;
m[13'd7578]=16'h0016;
m[13'd7579]=16'h090c;
m[13'd7580]=16'h000a;
m[13'd7581]=16'h090d;
m[13'd7582]=16'h0007;
m[13'd7583]=16'h000b;
m[13'd7584]=16'h000a;
m[13'd7585]=16'h410b;
m[13'd7586]=16'h0095;
m[13'd7587]=16'h000a;
m[13'd7588]=16'h0009;
m[13'd7589]=16'h5009;
m[13'd7590]=16'h007c;
m[13'd7591]=16'h0601;
m[13'd7592]=16'h0009;
m[13'd7593]=16'h6c00;
m[13'd7594]=16'h0018;
m[13'd7595]=16'h4104;
m[13'd7596]=16'h0025;
m[13'd7597]=16'h4004;
m[13'd7598]=16'h004e;
m[13'd7599]=16'h0003;
m[13'd7600]=16'h0009;
m[13'd7601]=16'hb002;
m[13'd7602]=16'h4a14;
m[13'd7603]=16'h810b;
m[13'd7604]=16'h002b;
m[13'd7605]=16'h3108;
m[13'd7606]=16'h0007;
m[13'd7607]=16'h0007;
m[13'd7608]=16'h0060;
m[13'd7609]=16'h000a;
m[13'd7610]=16'h0009;
m[13'd7611]=16'h6009;
m[13'd7612]=16'h0074;
m[13'd7613]=16'h0601;
m[13'd7614]=16'h0009;
m[13'd7615]=16'h6c00;
m[13'd7616]=16'h0018;
m[13'd7617]=16'h4104;
m[13'd7618]=16'h0025;
m[13'd7619]=16'h4004;
m[13'd7620]=16'h004e;
m[13'd7621]=16'h0003;
m[13'd7622]=16'h0009;
m[13'd7623]=16'hc002;
m[13'd7624]=16'h4b1e;
m[13'd7625]=16'h110b;
m[13'd7626]=16'h002b;
m[13'd7627]=16'h1108;
m[13'd7628]=16'h0007;
m[13'd7629]=16'h0007;
m[13'd7630]=16'h0060;
m[13'd7631]=16'h000a;
m[13'd7632]=16'h0009;
m[13'd7633]=16'h7009;
m[13'd7634]=16'h0074;
m[13'd7635]=16'h0601;
m[13'd7636]=16'h0009;
m[13'd7637]=16'h6c00;
m[13'd7638]=16'h0018;
m[13'd7639]=16'h4104;
m[13'd7640]=16'h0025;
m[13'd7641]=16'h4004;
m[13'd7642]=16'h004e;
m[13'd7643]=16'h0003;
m[13'd7644]=16'h0009;
m[13'd7645]=16'hd002;
m[13'd7646]=16'h4b1b;
m[13'd7647]=16'h800b;
m[13'd7648]=16'h002b;
m[13'd7649]=16'h0808;
m[13'd7650]=16'h0007;
m[13'd7651]=16'h0007;
m[13'd7652]=16'h0060;
m[13'd7653]=16'h000a;
m[13'd7654]=16'h0009;
m[13'd7655]=16'h8009;
m[13'd7656]=16'h0074;
m[13'd7657]=16'h0601;
m[13'd7658]=16'h0009;
m[13'd7659]=16'h6c00;
m[13'd7660]=16'h0018;
m[13'd7661]=16'h4104;
m[13'd7662]=16'h0025;
m[13'd7663]=16'h4004;
m[13'd7664]=16'h004e;
m[13'd7665]=16'h0003;
m[13'd7666]=16'h0009;
m[13'd7667]=16'he002;
m[13'd7668]=16'h4b1b;
m[13'd7669]=16'h400b;
m[13'd7670]=16'h002b;
m[13'd7671]=16'h1608;
m[13'd7672]=16'h0007;
m[13'd7673]=16'h0007;
m[13'd7674]=16'h0060;
m[13'd7675]=16'h000a;
m[13'd7676]=16'h0009;
m[13'd7677]=16'h9009;
m[13'd7678]=16'h0074;
m[13'd7679]=16'h0601;
m[13'd7680]=16'h0009;
m[13'd7681]=16'h6c00;
m[13'd7682]=16'h0018;
m[13'd7683]=16'h4104;
m[13'd7684]=16'h0025;
m[13'd7685]=16'h4004;
m[13'd7686]=16'h004e;
m[13'd7687]=16'h0003;
m[13'd7688]=16'h0009;
m[13'd7689]=16'hf002;
m[13'd7690]=16'h4b1e;
m[13'd7691]=16'h800b;
m[13'd7692]=16'h002b;
m[13'd7693]=16'h0508;
m[13'd7694]=16'h0007;
m[13'd7695]=16'h0007;
m[13'd7696]=16'h0060;
m[13'd7697]=16'h000a;
m[13'd7698]=16'h0009;
m[13'd7699]=16'ha009;
m[13'd7700]=16'h0074;
m[13'd7701]=16'h0601;
m[13'd7702]=16'h0009;
m[13'd7703]=16'h6c00;
m[13'd7704]=16'h0018;
m[13'd7705]=16'h4104;
m[13'd7706]=16'h0025;
m[13'd7707]=16'h4004;
m[13'd7708]=16'h004e;
m[13'd7709]=16'h0103;
m[13'd7710]=16'h0009;
m[13'd7711]=16'h0002;
m[13'd7712]=16'h4b2b;
m[13'd7713]=16'h800b;
m[13'd7714]=16'h002b;
m[13'd7715]=16'h0408;
m[13'd7716]=16'h0007;
m[13'd7717]=16'h0007;
m[13'd7718]=16'h0025;
m[13'd7719]=16'h400b;
m[13'd7720]=16'h004e;
m[13'd7721]=16'h000a;
m[13'd7722]=16'h0009;
m[13'd7723]=16'hb009;
m[13'd7724]=16'h0110;
m[13'd7725]=16'h0501;
m[13'd7726]=16'h0009;
m[13'd7727]=16'hb900;
m[13'd7728]=16'h001b;
m[13'd7729]=16'h4002;
m[13'd7730]=16'h0010;
m[13'd7731]=16'h0003;
m[13'd7732]=16'h0016;
m[13'd7733]=16'h0905;
m[13'd7734]=16'h000a;
m[13'd7735]=16'h0906;
m[13'd7736]=16'h0007;
m[13'd7737]=16'h0004;
m[13'd7738]=16'h000a;
m[13'd7739]=16'h4104;
m[13'd7740]=16'h008d;
m[13'd7741]=16'h0003;
m[13'd7742]=16'h0009;
m[13'd7743]=16'h5002;
m[13'd7744]=16'h49ff;
m[13'd7745]=16'h800b;
m[13'd7746]=16'h002b;
m[13'd7747]=16'h0308;
m[13'd7748]=16'h0007;
m[13'd7749]=16'h0007;
m[13'd7750]=16'h0025;
m[13'd7751]=16'h400b;
m[13'd7752]=16'h004e;
m[13'd7753]=16'h000a;
m[13'd7754]=16'h0009;
m[13'd7755]=16'hc009;
m[13'd7756]=16'h0055;
m[13'd7757]=16'h4801;
m[13'd7758]=16'h0007;
m[13'd7759]=16'h0000;
m[13'd7760]=16'h000e;
m[13'd7761]=16'h8104;
m[13'd7762]=16'h0058;
m[13'd7763]=16'h0003;
m[13'd7764]=16'h0009;
m[13'd7765]=16'h6002;
m[13'd7766]=16'h4b4e;
m[13'd7767]=16'h800b;
m[13'd7768]=16'h002b;
m[13'd7769]=16'h0308;
m[13'd7770]=16'h0007;
m[13'd7771]=16'h0007;
m[13'd7772]=16'h0025;
m[13'd7773]=16'h400b;
m[13'd7774]=16'h004e;
m[13'd7775]=16'h000a;
m[13'd7776]=16'h0009;
m[13'd7777]=16'hd009;
m[13'd7778]=16'h0074;
m[13'd7779]=16'h0501;
m[13'd7780]=16'h0009;
m[13'd7781]=16'hb900;
m[13'd7782]=16'h0018;
m[13'd7783]=16'h4104;
m[13'd7784]=16'h0058;
m[13'd7785]=16'h0003;
m[13'd7786]=16'h0009;
m[13'd7787]=16'h7002;
m[13'd7788]=16'h4b24;
m[13'd7789]=16'h100b;
m[13'd7790]=16'h002b;
m[13'd7791]=16'h1208;
m[13'd7792]=16'h0007;
m[13'd7793]=16'h0007;
m[13'd7794]=16'h0025;
m[13'd7795]=16'h400b;
m[13'd7796]=16'h004e;
m[13'd7797]=16'h000a;
m[13'd7798]=16'h0009;
m[13'd7799]=16'he009;
m[13'd7800]=16'h0074;
m[13'd7801]=16'h0501;
m[13'd7802]=16'h0009;
m[13'd7803]=16'hb900;
m[13'd7804]=16'h0018;
m[13'd7805]=16'h4104;
m[13'd7806]=16'h0058;
m[13'd7807]=16'h0003;
m[13'd7808]=16'h0009;
m[13'd7809]=16'h8002;
m[13'd7810]=16'h4b24;
m[13'd7811]=16'h100b;
m[13'd7812]=16'h002b;
m[13'd7813]=16'h1208;
m[13'd7814]=16'h0007;
m[13'd7815]=16'h0007;
m[13'd7816]=16'h0025;
m[13'd7817]=16'h400b;
m[13'd7818]=16'h004e;
m[13'd7819]=16'h000a;
m[13'd7820]=16'h0009;
m[13'd7821]=16'hf009;
m[13'd7822]=16'h0074;
m[13'd7823]=16'h0501;
m[13'd7824]=16'h0009;
m[13'd7825]=16'hb900;
m[13'd7826]=16'h0018;
m[13'd7827]=16'h4104;
m[13'd7828]=16'h0058;
m[13'd7829]=16'h0003;
m[13'd7830]=16'h0009;
m[13'd7831]=16'h9002;
m[13'd7832]=16'h4b24;
m[13'd7833]=16'h100b;
m[13'd7834]=16'h002b;
m[13'd7835]=16'h1108;
m[13'd7836]=16'h0007;
m[13'd7837]=16'h0007;
m[13'd7838]=16'h0025;
m[13'd7839]=16'h400b;
m[13'd7840]=16'h004e;
m[13'd7841]=16'h010a;
m[13'd7842]=16'h0009;
m[13'd7843]=16'h0009;
m[13'd7844]=16'h0074;
m[13'd7845]=16'h0501;
m[13'd7846]=16'h0009;
m[13'd7847]=16'hb900;
m[13'd7848]=16'h0018;
m[13'd7849]=16'h4104;
m[13'd7850]=16'h0058;
m[13'd7851]=16'h0003;
m[13'd7852]=16'h0009;
m[13'd7853]=16'ha002;
m[13'd7854]=16'h4bae;
m[13'd7855]=16'h0608;
m[13'd7856]=16'h0009;
m[13'd7857]=16'h6c07;
m[13'd7858]=16'h001b;
m[13'd7859]=16'h4009;
m[13'd7860]=16'h0010;
m[13'd7861]=16'h000a;
m[13'd7862]=16'h0016;
m[13'd7863]=16'h090c;
m[13'd7864]=16'h000a;
m[13'd7865]=16'h090d;
m[13'd7866]=16'h0007;
m[13'd7867]=16'h000b;
m[13'd7868]=16'h000a;
m[13'd7869]=16'h410b;
m[13'd7870]=16'h0095;
m[13'd7871]=16'h000a;
m[13'd7872]=16'h0009;
m[13'd7873]=16'h5009;
m[13'd7874]=16'h0103;
m[13'd7875]=16'h0601;
m[13'd7876]=16'h0009;
m[13'd7877]=16'h6c00;
m[13'd7878]=16'h001b;
m[13'd7879]=16'h4002;
m[13'd7880]=16'h0010;
m[13'd7881]=16'h0003;
m[13'd7882]=16'h0016;
m[13'd7883]=16'h0905;
m[13'd7884]=16'h000a;
m[13'd7885]=16'h0906;
m[13'd7886]=16'h0007;
m[13'd7887]=16'h0004;
m[13'd7888]=16'h000a;
m[13'd7889]=16'h4104;
m[13'd7890]=16'h008d;
m[13'd7891]=16'h0003;
m[13'd7892]=16'h0009;
m[13'd7893]=16'h5002;
m[13'd7894]=16'h4978;
m[13'd7895]=16'h000a;
m[13'd7896]=16'h0009;
m[13'd7897]=16'h6009;
m[13'd7898]=16'h0055;
m[13'd7899]=16'h4801;
m[13'd7900]=16'h0007;
m[13'd7901]=16'h0000;
m[13'd7902]=16'h000e;
m[13'd7903]=16'h8104;
m[13'd7904]=16'h0058;
m[13'd7905]=16'h0003;
m[13'd7906]=16'h0009;
m[13'd7907]=16'h6002;
m[13'd7908]=16'h4bf3;
m[13'd7909]=16'h000a;
m[13'd7910]=16'h0009;
m[13'd7911]=16'h7009;
m[13'd7912]=16'h0074;
m[13'd7913]=16'h0601;
m[13'd7914]=16'h0009;
m[13'd7915]=16'h6c00;
m[13'd7916]=16'h0018;
m[13'd7917]=16'h4104;
m[13'd7918]=16'h0058;
m[13'd7919]=16'h0003;
m[13'd7920]=16'h0009;
m[13'd7921]=16'h7002;
m[13'd7922]=16'h4bc9;
m[13'd7923]=16'h000a;
m[13'd7924]=16'h0009;
m[13'd7925]=16'h8009;
m[13'd7926]=16'h0074;
m[13'd7927]=16'h0601;
m[13'd7928]=16'h0009;
m[13'd7929]=16'h6c00;
m[13'd7930]=16'h0018;
m[13'd7931]=16'h4104;
m[13'd7932]=16'h0058;
m[13'd7933]=16'h0003;
m[13'd7934]=16'h0009;
m[13'd7935]=16'h8002;
m[13'd7936]=16'h4bc9;
m[13'd7937]=16'h000a;
m[13'd7938]=16'h0009;
m[13'd7939]=16'h9009;
m[13'd7940]=16'h0074;
m[13'd7941]=16'h0601;
m[13'd7942]=16'h0009;
m[13'd7943]=16'h6c00;
m[13'd7944]=16'h0018;
m[13'd7945]=16'h4104;
m[13'd7946]=16'h0058;
m[13'd7947]=16'h0003;
m[13'd7948]=16'h0009;
m[13'd7949]=16'h9002;
m[13'd7950]=16'h4bc9;
m[13'd7951]=16'h000a;
m[13'd7952]=16'h0009;
m[13'd7953]=16'ha009;
m[13'd7954]=16'h0074;
m[13'd7955]=16'h0601;
m[13'd7956]=16'h0009;
m[13'd7957]=16'h6c00;
m[13'd7958]=16'h0018;
m[13'd7959]=16'h4104;
m[13'd7960]=16'h0058;
m[13'd7961]=16'h0003;
m[13'd7962]=16'h0009;
m[13'd7963]=16'ha002;
m[13'd7964]=16'h4b9e;
m[13'd7965]=16'h400b;
m[13'd7966]=16'h004e;
m[13'd7967]=16'h000a;
m[13'd7968]=16'h0009;
m[13'd7969]=16'hb009;
m[13'd7970]=16'h0103;
m[13'd7971]=16'h0601;
m[13'd7972]=16'h0009;
m[13'd7973]=16'hce00;
m[13'd7974]=16'h001b;
m[13'd7975]=16'h4002;
m[13'd7976]=16'h0010;
m[13'd7977]=16'h0003;
m[13'd7978]=16'h0016;
m[13'd7979]=16'h0905;
m[13'd7980]=16'h000a;
m[13'd7981]=16'h0906;
m[13'd7982]=16'h0007;
m[13'd7983]=16'h0004;
m[13'd7984]=16'h000a;
m[13'd7985]=16'h4104;
m[13'd7986]=16'h008d;
m[13'd7987]=16'h0003;
m[13'd7988]=16'h0009;
m[13'd7989]=16'h5002;
m[13'd7990]=16'h4a63;
m[13'd7991]=16'h400b;
m[13'd7992]=16'h004e;
m[13'd7993]=16'h000a;
m[13'd7994]=16'h0009;
m[13'd7995]=16'hc009;
m[13'd7996]=16'h0055;
m[13'd7997]=16'h4801;
m[13'd7998]=16'h0007;
m[13'd7999]=16'h0000;
m[13'd8000]=16'h000e;
m[13'd8001]=16'h8104;
m[13'd8002]=16'h0058;
m[13'd8003]=16'h0003;
m[13'd8004]=16'h0009;
m[13'd8005]=16'h6002;
m[13'd8006]=16'h4ba6;
m[13'd8007]=16'h400b;
m[13'd8008]=16'h004e;
m[13'd8009]=16'h000a;
m[13'd8010]=16'h0009;
m[13'd8011]=16'hd009;
m[13'd8012]=16'h0074;
m[13'd8013]=16'h0601;
m[13'd8014]=16'h0009;
m[13'd8015]=16'hce00;
m[13'd8016]=16'h0018;
m[13'd8017]=16'h4104;
m[13'd8018]=16'h0058;
m[13'd8019]=16'h0003;
m[13'd8020]=16'h0009;
m[13'd8021]=16'h7002;
m[13'd8022]=16'h4b7c;
m[13'd8023]=16'h400b;
m[13'd8024]=16'h004e;
m[13'd8025]=16'h000a;
m[13'd8026]=16'h0009;
m[13'd8027]=16'he009;
m[13'd8028]=16'h0074;
m[13'd8029]=16'h0601;
m[13'd8030]=16'h0009;
m[13'd8031]=16'hce00;
m[13'd8032]=16'h0018;
m[13'd8033]=16'h4104;
m[13'd8034]=16'h0058;
m[13'd8035]=16'h0003;
m[13'd8036]=16'h0009;
m[13'd8037]=16'h8002;
m[13'd8038]=16'h4b79;
m[13'd8039]=16'h400b;
m[13'd8040]=16'h004e;
m[13'd8041]=16'h000a;
m[13'd8042]=16'h0009;
m[13'd8043]=16'hf009;
m[13'd8044]=16'h0074;
m[13'd8045]=16'h0601;
m[13'd8046]=16'h0009;
m[13'd8047]=16'hce00;
m[13'd8048]=16'h0018;
m[13'd8049]=16'h4104;
m[13'd8050]=16'h0058;
m[13'd8051]=16'h0003;
m[13'd8052]=16'h0009;
m[13'd8053]=16'h9002;
m[13'd8054]=16'h4b7c;
m[13'd8055]=16'h400b;
m[13'd8056]=16'h004e;
m[13'd8057]=16'h010a;
m[13'd8058]=16'h0009;
m[13'd8059]=16'h0009;
m[13'd8060]=16'h0074;
m[13'd8061]=16'h0601;
m[13'd8062]=16'h0009;
m[13'd8063]=16'hce00;
m[13'd8064]=16'h0018;
m[13'd8065]=16'h4104;
m[13'd8066]=16'h0058;
m[13'd8067]=16'h0003;
m[13'd8068]=16'h0009;
m[13'd8069]=16'ha002;
m[13'd8070]=16'h4c1a;
m[13'd8071]=16'h000f;
m[13'd8072]=16'h0009;
m[13'd8073]=16'h000e;
m[13'd8074]=16'h001b;
m[13'd8075]=16'h0010;
m[13'd8076]=16'h0010;
m[13'd8077]=16'h0011;
m[13'd8078]=16'h0015;
m[13'd8079]=16'h0013;
m[13'd8080]=16'h0009;
m[13'd8081]=16'h0014;
m[13'd8082]=16'h0007;
m[13'd8083]=16'h0012;
m[13'd8084]=16'h0009;
m[13'd8085]=16'h4012;
m[13'd8086]=16'h01e0;
m[13'd8087]=16'h0708;
m[13'd8088]=16'h0009;
m[13'd8089]=16'h3507;
m[13'd8090]=16'h001b;
m[13'd8091]=16'h4009;
m[13'd8092]=16'h0010;
m[13'd8093]=16'h000a;
m[13'd8094]=16'h0016;
m[13'd8095]=16'h090c;

end

endmodule
